��Ȏظ ���1����\|                               BOOTLOADER ERROR, STAGE 0
                 ��|� ���U�|�A��� ��U��� 1�� ~f�   �� f� ~  fg�Ff�|fg�Ff�|fg�F f�|fg�F(f� |fg�F,f�$|f�|f�(|f�$|f�&|f(|f�,|1�� ~f�,|�k f� ~  fg�Fkf�&|f(|f��fg�Fof1�f�6|f��f�1�� ��8 f��|��1Ҋ|f��}fSR� �  �0|� 1���`��< t����a�f`�L|��D �D �\�|f�Df�D    �|�B�rfa�fa뱐��������������������������������������������������������  ����������������                                                U�KINGUIO_                         �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ������������������������      	   
                  ����                                                 !   "   #   $   %   &   '   (   )   *   +   ,   -   ������������1   2   3   4   5   6   7   8   9   :   ;   <   =   ����?   @   A   B   C   D   E   F   G   H   I   J   ����L   M   N   O   P   Q   R   S   T   U   V   W   ����Y   Z   [   \   ]   ^   _   `   a   b   c   d   e   ����g   h   i   j   k   l   m   n   o   p   q   r   s   ����u   v   w   x   y   z   {   |   }   ~      �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �������������������������   �   �   �   �   �   �   �   �   �   �   �����   �   �   �   �   �   �   �   �   �   �   �����   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �����   �   �   �   �   �   �   �   �   �   �   �   �   ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                stage1.bin                                                                                       �            ^
               bin                                                                                              �@                           system                                                                                           �@                           user                                                                                             �@                           stage2.bin                                                                                       �            d7             kernel.bin                                                                                       �            `�             ap.bin                                                                                           �         .                  README.md                                                                                        �         /   .               term.bin                                                                                         �         0   h�             shell.bin                                                                                        �         >   �� 	            launcher.bin                                                                                     �         K   0� 
            explore.bin                                                                                      �         X   ��             editor.bin                                                                                       �         f   ��             logo.bmp                                                                                         �         t   ��             folder.bmp                                                                                       �         �   �              console.bmp                                                                                      �         �   �              edit.bmp                                                                                         �         �   �              file.bmp                                                                                         �         �   �              text.bmp                                                                                         �         �   �              test.bin                                                                                         �         �   �v             cat.bin                                                                                          �         �    w             lua.bin                                                                                          �         �   @             nanojpeg.bin                                                                                     �         �   ��             test.lua                                                                                         �         �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��  BOOTLOADER ERROR, STAGE 1 Sirius Boot Manager Version 2.0
 BM-SHELL:/>  install system boot                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               stage2.bin                                                                                       kernel.bin                                                                                       ap.bin                                                                                           `��< t����a�1�����READ ERROR
 f`�h���D �D �\�|f�Df�D    �b��B�rfa�a�����WRITHE ERROR
 f`�x���D �D �\�|f�Df�D    �g�� �C�rfa�a�0��[���|�f�������1�� ~f�   �c�f� ~  fg�Ff���fg�Ff���fg�F f���fg�F,f���f���f���f���f�&��f��f���1����f���f�����1ҋ6���>���@ 1Ɋ�%8�u
AFG��`t"��1Ɂ �>���6��փ� t��1��Ҹ Ë6���f�Dkf������f���f�&��f��f����>�������������&��� �)Á� 9��t���  ����  ��� f�   f�&��f1�f�6��f��1�� ~�M�f1�f���f�   f��f1�f��f���f�� �� ~�f�f���f���t�X�1��BIOSes Extensions Parameters not present
 BIOSes Get Device Parameters Error
 BIOSes Enhanced disk device not suport (EDD)
 �A�b���U�s��U�t���=�� u�5��2� �J �H�b���� t���VW� @��1��J ��_^����`��5 ����/ ���d�! �`���! ���d� ���`� ���d�
 �a��d�t���d�u��VESA VBE ERROR
     �� ��O�1��޾ � @��1�� ������ ��O�� ��8��t�	�����g����>1ۋ�������t#� ��O�� ��8��t�	��9��}/���π>� u�>� t�� �� 1�뱀.�1���e1��޾��� @�ǿ � ��f1ۋ��� @�2 ��Ou:�f1�W� O� f�VBE2�_�f1��  ��W�O����_�f1�W�O�_þ����1���`�O�1�1Ҏ¿ �a�        ��   �� ��   �� ��   �  ��   �  ' F�  VW��$8�u	�� tGF��_^þ��C��A��=�� QP�  �  �����XY� �2�<t�G���
����� �]����� t� �N����� t��Q� @1�� f�    ���H�f����Y����Ȏ؎�� ���1�����b�f�c��g���g���=���f�c�    ���  ����>����� ��� ���  ���  �,��� t���m�1������  �r��>����� ��� @���  ���  ����� t���4�1������  ���>����� ��� P���  ���  ���� t�����1����N��2���p��pf�n�  fg �f��"�f1Ҋb�f�c�f1ɋ��f�6�   1�`�=2�  �< t��f���a� � �   �؎�����м  	 �    �  SQRT�P��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ELF                4   �4     4    (              �   �            �   �  �     �           �   �  �               Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �    � p �    �<p �@p �z �   �U��D$�8  f� f��f��f��f��f�Љ�]�U��D$��]�U��D$�T$�\$��]��      ��H1ɉ�M1�M1�M1�M1�M1�M1�M1�M1�H1�H� p     H1�f��f��f��f��f���H1ۉÉ�S�����������L$����q�U��SQ��`��  ���  ��h   ��  ���c  ����<���P�l  �����E�P�uZ  �����E�P��m���P�G  ������<���P�5  ����Dp � �H��Dp � �PD��Dp � �@@QRP��q���P�  ������<���P��  ����������P��  ����  �  ����<���P��  ���    �怃���<���P�  ���O:  ����<���P�  ����jj �K"  ����<p � ������@p �  ����<���P�[  ����������P�I  ����z � ����   ��������P������P�  ���E�}� u��������P�  ������jj �u��  �����u��  ���E����u��  ���E��u�Pjh  @ �  �����u��`  ���!��z � ����Ph   h  @ �  ������<���P�y
  �����E�P�E�Ph  ��GY  ���E�%    ��u��������P��	  ������������P��	  ���Z  ����<���P�
  ���7`  �E���u�h @ ��  ����e�Y[]�a����U����b�  ^�  �M���Q����������)ЉE��怃m��}� u�������U���$�   �  �� p �U��]���U����  �  �� p �
�U��� p �
�� p � +E]���U���ҋ  ��  �]���U��S��趋  �ö�  �} u�E�E�E�P�U�� 0�E��  ��   �E�E�U�EЉE��/�E���E��m��}�	~�7   ��0   �U�Ѓm��E��E�;EwɋU�E��  �E�E��E�    �'�E�� <0u�E�����u��u��  ����E��E�;E|ыE�E���u��!  ���E�   +E�M�U�ʃ�Pj R�  ���]�����U��� 贊  ��  �E�E��E�E��E�    �}� y)�E��P�U�� -�}�   �u�E�����E���E��؉E��E��E��M��gfff����������)�����)��ʉЍH0�E��P�U��ʈ�M��gfff����������)ЉE��}� u��}� t�E�� ���E���E��P��U��  �)�E�� �E�E��P�U��U����E��P��U��U��E�;E�wϋE����U���訉  ��  �E�E�E�E��E�E���E��P�U��U��m��}� u�E����U����b�  ^�  �E�E��E�E��E�E���U�B�E�E��H�M����E��P��U���u܋E����U�����  �  �E�E�E�E��E�E���U��B�E��E��H�M����E�� ��uߋE��  �E�����U���轈  ��  �E�E���E��E�� ��u�E�+E����U��S��膈  �Æ�  ��jd�i�������Dp ���Dp � ��jdj P�������E�  �E�  �E������Dp � �҉�E������Dp � �҉P�E������Dp � �҉P�E������Dp � �҉P�E������Dp � �҉P��Dp ���Dp � �R�P��Dp � �@    ��Dp � �U��R(�P �E�����Dp � �҉P��h  � �l���������Dp � �P(��Dp ���Dp � �R �P0��Dp � �@8    ��Dp � �@<    ��Dp ���Dp � �R�P@��Dp ���Dp � �R�PD��Dp ���Dp � �R�P��Dp � �@P   ��Dp � �@T   ��Dp � �@X��� ��Dp � �@\    ��Dp � �� � �P`��]�����U��蘆  ��  ��Dp ��J�U�ʋU�����Dp � �@0ЉE��]���U����T�  P�  �U�U���Dp ��J�U9�v8��Dp ��R��u)��Dp � �P�E�ЋEЍ�    �E�E�������U��S����  ��  ��Dp ��J@��Dp ��RD����Dp ��R������Dp �	�I(����Dp �	�I0��RSQ���'�������]�����U��S���{�  ��{�  ��Dp � �P@��Dp � �@D����Dp � �@������Dp ��R0��Pj R��������Dp � �@L    ��Dp ��@L�BH��]�����U�����  ��  f�E�  �E�@�E��E�    �of�E� �E�@�E�E�Ѝ �E��� f�E�E� ���E��2�E�f#E�f��t�U�E�M�E���uRP�������f�e��m��}� yȃE��E�@9E�|�������U��WVS���R�  ��R�  �}
u(��Dp � �@H    ��Dp � �PL���PL�E�  �}�E�   ��Dp � �PL��Dp � �@T����Dp � �@D��9�r��Dp � �@L    ��Dp � �PH��Dp � �@P����Dp � �@@9�r ��Dp � �@H    ��Dp � �PL���PL��Dp � �pP��Dp � �@(�E���Dp � �HX��Dp � �PL��Dp � �@T����Dp � �PH��Dp � �@P��V�u�Q�uWP��������Dp � �PH���PH�E�e�[^_]���U��S�����  ��  ���u���������]�����U��S���΂  ����  �} t>�E�    ��U�E�� ����P�������E����u��������U�9�w����]�����U��S��  �k�  ��k�  ��h   j ������P�������E�E�E���u�P������P�h  ���E���������P�=������E��]�����U��S����   �  �U���u�    ����u�u���J  ���E�E�]�����U��S�����  ��  ���u���K  ���]�����U��蚁  ��  �} t1�E�@"    �E�P"�E�P�Ef�   �E�@���E�P��]���U���O�  K�  �}tL�}g�} t�}t�Y�U�E�P�U�E�P"�E�E�P�EE�P�E�P"�EE�P"�!�E��&  �E)E�P�E�P�E�P"��E�@�U�J�    ��ЉEf��    ]���U��觀  ��  �} u�    ��E�@]���U��S��聀  ��y�  �E�P�E��&  9�r
������   �E�@����u:�E�@���E�P�E�@�U�Z�    ��E���u��u���J  ���E�H�E� ���ӋUf����E�P�E�@� ���E��E� �ЋE�@9�r�E�@���E�P�Ef�   �E�@�P�E�P�E��]�����U����  ��  �} u�    �g�E�    �E�E��E�    �:���u��������E�}��u�E�    �u�-�E�P�U�U��E��E��E�E9E�r��E�    �u����U����  �  �E�E��E�E���U��B�E��E��H�M����E�� ��uߋE�����U��S��$  �~  �õ�  �E�E�f�E�  �E� �E�    �  �U��E�� ����%�V  �E��U��E�� ����X�� �  ��������>���E�E��� �E��E�E��E�P�u��������E���   �E�E�@��E��u��u���������E���   �E�E�@��E��������P�u��!�������������P�u��������E��   �E�E��� �E��E��������RP���������������P�u��x������E��X�E�E�@��E�E��j������RP��������������P�u��9������E���������P�u��������E���$�U��E�� �E����E�P�u���������E���E��U��E�� ���X����U�E)Ћ]�����U��WVS��(��|  ʼ  �E�M�u �uЋ}$�}̋}(�u,�]0�U4�E��ȈE��EЈE��ËE���E����E܉؈E؉ЈEԋE��    �EЋU������� 	وf�����P�� 	ʈP�E��    �EЋU�����H�� 	وHf�����P�� 	ʈP�E�����E��    �EЉʈP�E��    �E��U����у��P���	ʈP�E��    �E��U���������P���	ʈP�E��    �E��U���������P��	ʈP�E��    �E��U�������P��	ʈP�E�����E��    �Eȃ������B���	ȈB�E��    �E��U����������P���	ʈP�E��    �E��U܃��������P���	ʈP�E��    �E��U؃��������P��	ʈP�E��    �E��Uԃ������P��	ʈP�E�����E��    �EЉʈP���([^_]���U��S���Lz  ��L�  ��jj ��xp P������j j j j j j j j j j j ��xp P�2�����0jjj j jj jj
j h�� j��xp P�
�����0jjj j jj jjj h�� j��xp P�������0��Hp f�  ��xp �    ��Hp �A�Q����Hp P��������]�����U��S���qy  ��q�  ��jj ��Tp P������j j j j j j j j j j j ��Tp P�W�����0j j jj jj jj
j j j��Tp P�2�����0j j jj jj jjj j j��Tp P������0��lp f�  ��Tp �    ��lp �A�Q���u�u��lp P��������]�����U��WVS���x  ��  �U�u�]�Mf�U���U�ڈU�ʈU�U��� p �Mf�]������ʃ� ��	������]�f�����\��� 	�\�� p �M�u��\��� 	�\��u��\��� 	�\�� p �M�D� �U����� p �M�ރ��\����	�\��U����� p �M�������\���	�\��U����� p �M�����\���	�\��U�������p �U�����\��� 	�\�f�����L��� 	وL����[^_]���U��S���/w  ��/�  ��h   j ���p P�`�������  ��  ���x f� ����p �    ���x �A�Q�����x P�$�������]�����U�����v  ��  �E�Uf�E��ЈE��U��E�jRh�   P�u�u������������U����|v  x�  �E�Uf�E��ЈE��U��E�jRh�   P�u�u���������f�`���D$4P�   f��f��f��f���  X��a��   �h    h    ����h    h   ����h    h   ����h    h   ����h    h   ����h    h   �s���h    h   �d���h    h   �U���h   �K���h    h	   �<���h
   �2���h   �(���h   ����h   ����h   �
���h    h   �����h    h   �����h   �����h    h   �����h    h   �����h    h   ����h    h   ����h    h   ����h    h   ����h    h   �y���h    h   �j���h    h   �[���h    h   �L���h    h   �=���h    h   �.���h    h   ����h    h   ����h    h    `���D$4P�   f��f��f��f���  X��a��   �h    h!   ����h    h"   ����h    h#   ����h    h$   ����h    h%   ����j j&�y���h    h'   �j���h    h(   �[���h    h)   �L���h    h*   �=���h    h+   �.���h    h,   ����h    h-   ����h    h.   ����h    h/   �������U��S���(s  ��(�  ���) j jPj �D�������* j jPj�/�������* j jPj�_������� * j jPj��������/* j jPj���������>* j jPj���������M* j jPj���������\* j jPj��������k* j jPj��������u* j jPj	���������* j jPj
�r��������* j jPj�]��������* j jPj�H��������* j jPj�3��������* j jPj���������* j jPj�	��������* j jPj����������* j jPj����������* j jPj����������* j jPj���������* j jPj$��������+ j jPj��������+ j jPj�v�������)+ j jPj�a�������8+ j jPj�L�������G+ j jPj�7�������V+ j jPj�"�������e+ j jPj��������t+ j jPj����������+ j jPj����������+ j jPj����������+ j jPj��������]�����U��S���lp  ��l�  �E���    ��P�u������}u* ЉE� ؉E� ��E��u��u��u�P���P����������U��S���p  ���  �D  ���+ j jPj �j��������+ j jPj!�U��������+ j jPj"�@�������, j jPj#�+�������, j jPj$��������), j jPj%��������8, j jPj&���������A, j jPj'���������P, j jPj(���������_, j jPj)��������n, j jPj*��������}, j jPj+���������, j jPj,�n��������, j jPj-�Y��������, j jPj.�D��������, j jPj/�/�������]�����U���n  ��  �]���U��S���n  ��  ���;X  ���[]���U����kn  g�  �m �} t�}�U����  �E��E��Ѓ}~�    ��   �    �    �����U����n  �  f�E����E�   ������Љ��E�!�f�E��}�!   ���E��U��E�!к!   ��"��   ���E��U��E�f����!к�   �����U����m  ��  f�E�  �E�   ����Љ��E�	�f�E��}�!   ���E��U��E�	к!   ��"��   ���E��U��E�f����	к�   �����U����m  �  �E��%  � �E��% � 	E��%   	E%�   	�   ���  ��  ���E��E�����U���l  ��  �E��%  � �E��% � 	E��%   	E%�   	�   ���  �E��  �]���U����cl  _�  �E��%  � �E��% � 	E��%   	E%�   	�   ���  ��  ���E��E�����U���l  �  �E��%  � �E��% � 	E��%   	E%�   	�   ���  �E��  �]���U��S��$�k  �å�  �E���������P���P�������E�    ��   �E�    ��   �E�    �   j�u��u��u���������E�}����   �E�    �X�E苄à  %��� �E���9�t�E��7�E苄ä  ��P��f���P�������u��u��u�i���P�h������	�}��   ~��}�   u!���u��u��u��u䍃x���P�6����� ���E��}��>����E��}��$����E��E�;E�����    �]�����U��� �mj  i�  �E������E�    �   �E�    �~�E�    �k�E���%  � �E���% � 	E���%   	�  ���  ��  ���E�E�E��E���9Eu�E���    �E�E�����.�E��}�~��E��}��x����E��}��   �^������������U��� �i  ��  �E������E�    �E�    �   �E�    �   �E�    �o�E���%  � �E���% � 	E���%   	�  ���  ��  ���E�E�E��E����E9�u�E���E�U���	ЉE�E��.�E��}�v��E��}��t����E��}��   �W������������U��� �h  ��  �E������E�    �   �E�    �   �E�    �y�E���%  � �E���% � 	E���%   	�  ���  ��  ���E�E�E��E���9Eu'�E�����9Eu�E���E�U���	ЉE�E��.�E��}�~��E��}��j����E��}��   �M������������U��� ��g  ڧ  �E������E�    �   �E�    �   �E�    �   �E���%  � �E���% � 	E���%   	�  ���  ��  ���E�E�E��E���9Eu5�E�����9Eu'�E�����9Eu�E���E�U���	ЉE�E��2�E��}��o����E��}��U����E��}��   �8������������U�����f  �  �Ef�E��    ����U�����f  ¦  �Ef�E��    ����U����f  ��  �E#E�E��E���!E��E�����U����~f  ��v�  �}v���z �U��Ѓ� �@�����E����z �U��Ѓ� �@�����E����z �U��Ѓ� �@�����E����z �U��Ѓ� �@�����E�������U�����e  �  ���z �U��Ѓ� �@�����E��E�������U���e  ��  ��u����������t�   ��u������%�   ��uӸ    ����U���he  d�  ��u�d���������t�   ��u�K�����%�   ��tӸ    ����U���!e  �  ��u����������t�   ��u����������uո    ����U����d  ؤ  ��u�����������t�   ��u����������tո    ����U��S�d  �Ò�  �u����������z �U��Ѓ� �@�P�E��u���������]�����U��S���Md  ��E�  ���z �U��Ѓ� �@���E��E��E��E��������z �]��ڃ� �R��E�%�   ���z �M��ʃ� �R�[]���U��W��c  ͣ  ���z �U��Ѓ� �P�E����E����fm�_]���U��V�c  ��  ���z �U��Ѓ� �P�E����E����fo�^]���U��S���Vc  ��V�  j �u�u�u�������E��  �U�f��E������  f�Pj�u�u�u��������E�E������  �P
�E������  �P���  �U�P	���  �@
<u���  �@<u���z �    �   ���  �@
<u.���  �@<u ���z �    ��������P������������  �@
<u���  �@<u���z �    �8��������P��������������P��������������P��������j�u�u�u��������E�E�����Pj�u�u�u������ ���  �@
<uc���  �@<uUj�u�u�u�������E�E�% �  ��t3j�u�u�u�e������E�E����Pj�u�u�u������ ���  �@
<��   ���  �@<��   j@�u�u�u�������E�E� � ���Pj@�u�u�u�L����� j�u�u�u��������E�E�% �  ��t3j�u�u�u�������E�E����Pj�u�u�u������� jH�u�u�u�������E�E����PjH�u�u�u������� j<�u�u�u�Q������E��  �U�P/�E������  �P0j�u�u�u���������  �Pj�u�u�u� ��������  �Pj�u�u�u����������  �Pj�u�u�u����������  �Pj �u�u�u���������  �Pj$�u�u�u���������  �P#�    �]�����U��S�_  ��  �U���z �]��ك�0�Q�U���z �]��ك��Q�U���z �]��ك� �Q�U���z �]��ك� �Q�U���z �]��ك� �Q�U ���z �M��ȃ�0��[]���U��S����^  ���  �u�������u���������z �U��Ѓ� �@�P�    ����z �U��Ѓ� �@�P�    ����z �U��Ѓ� �@�P�    ����z �U��Ѓ� �@�P�    ����z �U��Ѓ��@������z �M��ʃ� �R����u�������u�]�����h�   �u�e������u�t������E�@B ��u�������%�   ��t�E��P��U���u����u��������E�}� u
�    �   ���z �U��Ѓ� �@�����E��E�E����z �U��Ѓ� �@�����E��E�E��}�u�}��u�   �>�}�iu�}�u�   �+�}� u�}� u�   ��}�<u�}��u�   ��    �]�����U��S����\  ����  �u����������/  ����t����>�����u�����P�D�������h   �u�u����������u����������u�g������E� f��y���  ��   ���z �U��Ѓ� ��E�   � ��%   ��t�0   ��   ���z �U��Ѓ��H���z �U��Ѓ��@    ���z �U��Ѓ��    �D  ���u��$���P�h�������h�   �u�4��������u�@��������u���������h   �u�u����������u����������u�\������E� f��y�   ����  ���z �U��Ѓ� ����z �U��Ѓ��@   ���z �U��Ѓ��@    ���z �U��Ѓ��    �[���u��7���P�����������u��H���P�h����������z �U��Ѓ� �     ���u��[���P�:�������    �]�����U��S���Z  �Ú�  �E�E��E�E����z �U��Ѓ��@��0��  ��0�m  ���J  ���\  �E�����z �U��Ѓ� �@�P���E������z �U��Ѓ� �@�P���E��U����������z �U��Ѓ� �@�P���E��U����������z �U��Ѓ� �@�P������z �U��Ѓ��@�����E��U���������	ȃ�@���z �M��ʃ� �R������z �U��Ѓ��P���x � 9��[  ���z �U��Ѓ� �P���x � 9��7  �u���������z �U��Ѓ��P���x ����z �U��Ѓ� �P���x ���  ���z �U��Ѓ� �@�P�    �E��U����������z �U��Ѓ� �@�P���E��U��1҉����z �U��Ѓ� �@�P���E��U��1��������z �U��Ѓ� �@�P������z �U��Ѓ� �@�P�E�E������z �U��Ѓ� �@�P���E��U����������z �U��Ѓ� �@�P���E��U����������z �U��Ѓ� �@�P������z �U��Ѓ��@����@���z �M��ʃ� �R������z �U��Ѓ��P���x � 9�t���z �U��Ѓ� �P���x � 9�t_�u����������z �U��Ѓ��P���x ����z �U��Ѓ� �P���x �����u������P�������������]�����U��S����V  ��ߖ  �E�E��E�E����z �U��Ѓ� � ���  ���  ��t
��t�  ������  �u��u��u�u����������z �U��Ѓ��@��t����   ��   ���z �U��Ѓ��@��t��0t�#��j �u���������j$�u�x���������u�Q��������u��������t������b���z �U��Ѓ�� ��P�u�u����������u���������u��������t���������������������    �]�����U��S���uU  ��u�  �E�E��E�E����z �U��Ѓ� � ���g  ���e  ��t
��t�W  ������R  �u��u��u�u�k��������z �U��Ѓ��@��t���  �  ���z �U��Ѓ��@��t��0t�#��j0�u� ��������j4�u����������u����������u��������t
������   ���z �U��Ѓ�� ��P�u�u���������z �U��Ѓ��@��t��0t�)��h�   �u���������h�   �u�v���������u�O��������u���������t���������������������    �]�����U��S���S  �ÿ�  ��������P�,�������h   j ���z P���������h   �t������E���h   �a��������  ��j��������E�}��u��������P����������E�����E������E�������QRP�������E�}� t�������P�{����������  �@������  �@��u��  ��    ���,p ����  �@������  �@��u��  ��    ��� p ����  �@������  �@��u�p  ��    ���4p ����  �@������  �@��u�v  ��    ���0p ����  �@�������$p ����  �@#�������8p ����z � ��t���'  �J  ����-���P�\�������$p � ���� p � ����,p � ��QRPj j jj ������ ��$p � ���� p � ����,p � ��QRPj jjj������� ��$p � ������0p � ����4p � ��QRPjj jj������ ��$p � ������0p � ����4p � ��QRPjjjj�u����� �E�    ����u��u���������E��}�~����x � �������x ����x ��<����>���P�:�������8p � ��P�#   �������P���P���������    �]�����U��S���qP  ��q�  ��h   �Q����������x ���h   �7��������x ��U���x ����x � ��P��
  ����]�����U���P  �  �E�@���E�P��E�@% @  ��u�E�@����E�P��E�@% �  ��u�]���U���O  ��  ��E�@% �  ��u�E�@���E�P�E�@���E�P�]���U��S���gO  ��g�  �u�E��������x ��E��E�@    �E� ��h   j P�w������E� ��   �E�P�E�@    �E�@��h   j P�C��������x � ��   ���x ����u��������]�����U��WVS��4�N  ��  �}�u�]�]��M$�](���U܉�U��U�f�UԋU�UȋU �Ủ�f�UЉڈU��E�    �U�U�U��@�U�U��'�U��J����J�U��J�ᏈJ�U܉у��U�����J��	وJ�U��B �U��M؈J�U��MĈJ���z �M��ʃ� ���t����   �  �EԉE�P�EȉE�P�EȋU������E�P�EȋU������E�P�E��@@�EȋU������E�P�EȋỦ�1҉E�P	�EȋỦ�1����E�P
�E�f���E�P�EЉE�P�E�f���E�P��   �UԉыU�J�U�f���ыU�J���z �U��Ѓ�� �E�E�E�P�E����E�P�E��@@�E�� ��E��@ �EȋU������E�P�EȋU������E�P�EȋU������E�P�EȉE�P�E��@ �E��@ �E��@ �EЉE�P	�E��@
 �E��@ ����4[^_]���U���DL  @�  �U�E���   �Eǀ�       �Eǀ�       �E%��? �E�с���? ���   ��  ��	ʉ��   �E���   f��?�f���   �E���   �ʀ���   �]���U��WVS���K  �®�  �}�u�]�M �E$�E܉��E����E�]�M��E܈E��E������E�˃�����	و���z �U��Ѓ� � ���E����������	ʈ�E���E���������	ʈ�E���E�������	ʈ�E���E�у��P���	ʈP�E����E����P���	ʈP�E�P����P�E�P����P�E�P���P�E(�Ef�P�E�U,�P�E�@��   �E�P�E�@    ���[^_]���U��WVS��<�OJ  ��O�  �U�E�UĈE��E�    �E�    �E�@�����E� �E�j jj j j j j�u�j �u�B�����(�E܋@�E؋E��@��������Pj �u��%��������x � ��h�  P�u��p������E؉EԋE�� '�E����Eԉу��P���	ʈP�E��P�ʀ�P�E��@��UċEԈP�E�   ����ЉE�P8�-�E�@ ����t��������P��������������   �E��E�@ %�   ��t	�}�?B ~��}�@B u��������P������������   �E�P8�E�   �����!Ѕ�t(�E�@%   @��t׃�������P�:�����������I��E܋@=   t��������P������������"���x ��E܋@�����E�ǉ���    �e�[^_]���U��S��$�MH  ��M�  �E�@(�E��E������E�E����E��E�    �E�    �E�    �}�t
�������  �}�t
�������  �E�@$=  �	  �E�   �E�   ���x Pj j��u�a������E����z �M��ʃ� ����x ���   ��%   ��t�0   ��   ���z �U��Ѓ��H���x �@b�����������z �M��ȃ��P�E����z �M��ʃ�����x �@x�����z �M��ʉB���z �U��ЋP���x �@z��������z �M��ȉP�  �E�@$=���   �E�   �E�   ���x Pj j��u�G������E����z �M��ʃ� ��E����z �M��ʃ�����z �U��Ѓ��@   ���z �U��Ѓ��@0   ���z �U����@    �g�E�@$=<�u�E�   �E�    �J�E�@$=i�u�E�   �E�    �-�E�    �E�    ���u�����P�Z�����������   �E􋄃�  ��P�u��7���P�0������E���z �M��ʃ�0�B���z �U��Ѓ�0�@���z �M��ʃ��B�E����z �M��ʃ�0�B���z �U��Ћ@   ������z �M��ȉP�    �]�����U����E  �  �U������U��U����z �P�E�    �B�E�����EЃ��uP�X������E�����EЃ��u�P�S������E��E�;E�|��    ����U��WVS��,�D  �È�  �E�EЋE�E����z �U��Ћ@��x
������  �E�    �E�    �E�@�����E� �E�j jj j j j j�u��u�u�[�����(�E܋@�E؋E��@��������Pj �u��>��������z �U��Ѓ�� �E�P����x � ��RP�u��s��������z �U��Ѓ� � ��t��tM�x���z �U��Ѓ��@��u(�E����j P�u��u�j j%j�u��u������0�7������  ���z �U��Ѓ��@��u
�������   �������   �E�   ����ЉE�P8��E�@ ����t
������   �E��E�@ %�   ��t	�}�?B ~́}�@B u������{�E�P8�E�   �����!Ѕ�t�E�@%   @��t׸�����K��E܋P���z �M��ȃ�� �E9�t�    �"���x ��E܋@�����E�ǉ���    �e�[^_]���U��WVS��,�5B  ��5�  �E�EЋE�E����z �U��Ћ@��x
������  �E�    �E�    �E�@�����E� �E�j jj j j jj�u��u�u������(�E܋@�E؋E��@��������Pj �u����������x � ���z �M��ʃ���U�����U�ǉ������z �U��Ѓ�� �E�P����x � ��RP�u�����������z �U��Ѓ� � ��t��tM�x���z �U��Ѓ��@��u(�E����j P�u��u�j j5j�u��u������0�7�������   ���z �U��Ѓ��@��u
�������   ������   �E�   ����ЉE�P8��E�@ ����t
������   �E��E�@ %�   ��t	�}�?B ~́}�@B u������^�E�P8�E�   �����!Ѕ�t�E�@%   @��t׸�����.��E܋P���z �M��ȃ�� �E9�t�    ��    �e�[^_]���U��WVS��<��?  ���  �E�E��E�EċE��E��E�    �E�    �E���EЋE�E��E�    �   ���z �U��Ѓ���E������EԋŰEԍ4�Eܺ    ���x �	�}�������VjRPQ�u������ �E��E����z �U��Ѓ�� ��    �E�ЉE؃}� t�E��^�E��E�9E��e����E���EЃ}� t<�ŰE؍4�Eܺ    ���x �	�]����ك�V�u�RPQ�u������ �E��E��e�[^_]���U��WVS��<�>  �Í~  �E�E��E�EċE��E��E�    �E�    �E���EЋE�E��E�    �   ���z �U��Ѓ���E������EԋŰEԍ4�Eܺ    ���x �	�}�������VjRPQ�u������ �E��E����z �U��Ѓ�� ��    �E�ЉE؃}� t�E��^�E��E�9E��e����E���EЃ}� t<�ŰE؍4�Eܺ    ���x �	�]����ك�V�u�RPQ�u�%����� �E��E��e�[^_]���U��WVS��,�I=  ��I}  �E�EЋE�EԋE�E����z � ��t
��tm�   �E�    �U���z �U��Ѓ���E��ЋE���E�Ɖ����EЋU�����QRPj�u������� ��t������@�E��E�9Ew��-���u��u�u��u��u������ ��t��������������    �e�[^_]���U��WVS��,�f<  ��f|  �E�EЋE�EԋE�E����z � ��t
��tm�   �E�    �U���z �U��Ѓ���E��ЋE���E�Ɖ����EЋU�����QRPj�u�f����� ��t������@�E��E�9Ew��-���u��u�u��u��u������ ��t��������������    �e�[^_]���U���  �;  �{  �E�E��E�E��������E��E�    �1�E�� ��u�U��E���  ��E��P�U��M��U��� ��E��}�_~��E�    �'�E��P�U���E�P�U�� 8�t�   ��E��}�_~Ӹ    ����U��S����:  ���z  �E�@�    �]����uRPjS���Y����� �]�����U��VS�� �:  �Ûz  �E�P�E�@ЉE��E�P,�E�@ �ЋE�ЉE��h    �S������E��h    j �u�蕰�����E�    �M�I �u�6���u�RPQV������� �E��E�    �)�E����E�Ѓ��uP�f������E�}� t�E��}�?~����E����E�Ѓ�h�   P�u�W��������u��ܭ�����    �e�[^]���U��VS��0�9  �Öy  ��hB  �v������E���hB  j �u�踯�����E��@    ��h    �D������U��B�E�Po�E���&  �E�P�E���*  �E�P �E���.  �E��E���:  ��h   �������U���>  �E�@k�E��h    �Ѭ�����E��E������E�    �E�    �{  ��h   褬�����U���>  �M���ʉ�E���>  �U���Ћ �E؃�h   j �u���������E�    �
  �E�@ �E�E�@��E�P�E�4�    �E��ʉ�E���6  �P�E���6  �E��    �E�p�Ⱥ    ���E�@E�@ЉEԋE�;E�tR�EԺ    �M�	���u�RPjQ�s����� �EЃ}� t#���u��ݫ�������u��  ���    �}�EԉE��E�@�����E��    ��U�E��    �E�Ћ �E�}��u	�E�������E��}��  ������}��t�E��}��  �x��������u��N������E��e�[^]���U��S��4�7  ��w  ��h   �������E��h   j �u��-�������jj �E�P�������E�   ��@p � ���EЃ��E�P�u��������E��}� t���u�贪�����    �i���uj �E�P�u����� P������ �E��}� t���u��x������    �-���E�P�u����� P�������E���u��G������E�]�����U��S���6  ��v  �E�@��P�������E�    �:�E��>  �U���Ћ ��t.�E��>  �U���Ћ ��P�ة�����E��}��  ~����E��>  ��P賩�������u襩�����E    �    �]�����U��WVS���a5  ��Yu  �E��6  �E9�v�} u������w�E��>  �E���  ��H���
��Ћ �E�E����%�  )Ѝ�    �E�Ћ �E��E�p�E�    �]��.  �}��:  ��VRPSW���g����� �e�[^_]���U��WVS���4  �t  �E�E��E��x�E��p�    ��ЋU�����E����  �    ��[^_]���U��WVS���X4  Tt  �E�E��E����E��E��P�U܋E��x�  ���ƋE��0�E���E܉��E����E؋E��H�M��E��x�E��p�  ���U܋U؉�E����U܉�E��� �E؋E��X$�]��E��x(�E��p,�  ���U܋U؉�E����U܉�    ��[^_]���U��VS�3  �s  �E��ƋE�0�E��[^]���U��WVS���a3  ]s  �E���E��E�P�U�E�x�E��ƋE�0�E���E���E� ��[^_]���U���3  s  �E��2���E��E��    ]���U�����2  �r  �E�    �E�    �E��2�E��U��E	E��E	E��E��U��M0�    ����U��S���2  �r  �U"ڃ�jx����������]�����U���k2  gr  �E"ؐ]���U���Q2  Mr   ��� "��]���U���42  0r   �   �"��]���U��WVS��L�2  ��r  ��(����E䋇,����E���h @ j �u����,������E�    �E�    ��   �U������U������E������    �Ȁ���E��ÉEԋMЋ]ԋU��ȃ������B��	��B�������B�� 	��B�������B�� 	��B�������B�� 	��B�����ƃ��B���	��B�؃������B��	��B�����������B���	ȈB�E��E�   �E��}��;  ������Dp � �@ �E��E�    ��   �U������U������E������    �Ȁ���E��ÉE̋Mȋ]̋U��ȃ������B��	��B�������B�� 	��B�������B�� 	��B�������B�� 	��B�����ƃ��B���	��B�؃������B��	��B�����������B���	ȈB�E��E�   �E��}��  ������h   j �u����������,����E��E�    ��   �U������U������E������    �Ȁ���E��ÉEċM��]ċU�ȃ������B��	��B�������B�� 	��B�������B�� 	��B�������B�� 	��B�����ƃ��B���	��B�؃������B��	��B�����������B���	ȈB�E�   �E��E��}�������$�����h   j P�����������$���������$���������(����E܋E�����$������    �Ȁ���E��ÉE��M��]��ȃ������F��	ЈF�������F�� 	ЈF�������F�� 	ЈF�������F�� 	ЈF�������F���	ЈF�؃������F��	ЈF���������F���	ЈF�� �����h   j P����������� ��������� ��������� ���������$����E܋E����� ����    �À���]��E��E��U��Ã������Y��	�Y�������Y�� 	�Y�������Y�� 	�Y�������Y�� 	�Y�����ރ��Y���	�Y�Ӄ������Y��	�Y���������A���	ЈA��X����� �����P�/�������j h   h�  ����������E�����h�  ����������Dp � �@0  ���e�[^_]���U��S���G,  ��Gl  �E�   �E�   ��h   j �u��n�������<p ��E���@p � �U������E���� �����E���� ��ЉE�E�P�E��E�� �   �E��$�    �E��(�  0 �E��,�  @ ��Dp � �U��@��jdPR�������E�]�����U���u+  qk  �   �    �   ��   �    �!   �(   ��   �   �!   �   ��   �   �!   �   ��   ��   �!   ��   ��   �]���U�����*  �j  �E�'  �} u)�怸d   ���E��E�����u<�E��P��U���u��-�}u'�怸d   ���E��E�����t�E��P��U���uې����U���y*  uj  j�n������E�d   �����U��S���J*  ��Jj  �E�E��j�9�������   �d   ��j�!������E��`   ]�����U��S����)  �i  ��j ����������`   ���E��E��]�����U�����)  �i  �����E��}��u�    ��}��u��������h�   �4�����������U��S���w)  ��wi  ���� �     ���� �     ���� �  ���� �     ���� �    ��j�3������    �d   ��j �������`   ���E��E��E��M���j��������`   �d   ��j��������E��`   ��j���������   �d   ��j��������h�   �B�����������h�   �-������v�����h�   �������a�����j�S��������� ����� � ��jj P荞�������� � �    ���� � �@   ��j���������]�����U��S����'  ���g  ���� � ��t���� �     �`   ���E��e  �d   ���E��E����  ���  �������;  ���  ���� ���&  ���� � �H���� �
����   ����   ��t
��t#��   �`   ���E��E������ ���   ���� � ������t#�`   ���E��E� ��������� ��   �`   ���E��U����� ��   ���� � ���� ��t������� ��������� ���`   ���E��U����� ����� � ��x���� � ����@��u�!   ���� �     ����� �     ���[]���U��S�[&  Wf  ��Dp ��R@��0�����Dp ��RD��4������� ������ �
���� �ى
���� ��Z���� �
���� �)ˉىJ���� �
���� ��I�J���� �
���� ��ɉJ���� ����y���� ��    �$���� ��
��0���9�~���� ���0����
���� ��R��y���� � �@    �&���� ��J��4���9�~���� ���4����B�[]���U��S���+%  'e  ��j ���������`   ���E��E��]�����U��S����$  �d  �U�U��j����������E��`   ]�����U����$  �d  �u����E��}��u�    ��}��u��������h�   ������������U��S���o$  kd  ��j���9�������]�����U��S���I$  ��Ad  ���  ��~
ǁ�      �`   ���E��E��E����  �P���  ���� �]���E���y�}��t�}��u$ǁ�      ��}�*t�}�6uǁ�     �J�E���xB�}�Et<���  ��t���  ��u�E����������  ��E����������  ��[]���U��S���`#  ��`c  ��� � ��h   j P菙������` � ��h   j P�t������� � � ��h   j P�Y�������� � ��h   j P�>�������� � ��h   j P�#�������` � ��h   j P�������� ` � ��h   j P��������]�����U����"  �b  ��` �
�U���` �
�� � �U���` ��E)E������U���I"  Eb  �E�@ ���E�P �E�@ ����u��]���U���"  b  �E�@ ����E�P �E�@ ����t��]���U����!  �a  �E�@ ���E�P �]���U���!  �a  �E�@ ���E�P �]���U���!  �a  �E�@ �� �E�P ��E�@ �� ��t�]���U���a!  ]a  �E�@ ��߉E�P �]���U��S���4!  ��4a  �u�
������E�@ ���E�P ��h�� 蘔�������jd艔�����E�@ ����u��������P�Y�������]�����U��S���   �þ`  j �u�u�u聳�����E�E����� � ��E������� � �Pj�u�u�u�L������E�E�% ������� � �P�� � �@����� ��    �]�����U��S���-   ��-`  ��������P蚝������` �     ��h �  j �� � P�@�������j jj��������E��}��u��������P�������������  �E��ЋE������M�����RPQ��������� � �H�� � �P�� � � QRP������P�������� � �@�E�������P�Ҝ�������u�����������u����������u��d������E�@ ��߉E�P �E��@8   ��� � �P(��� � ���P(��h   �K�������� ���h   �3�������� ���h   ��������` ���h   �������� � ���h   ���������� ���h   ���������� ���h   ��������` ���h   �������� ` ���� � �    ��� � �@    ��� � �@    ��� � �@    ��� � �@   ��� � �@    ��� � �@    �E�    ���� � ������ p �U���E��}��  ~���� � �@0    ��� � �� p �P4��� � �@,    �E��@8    ��� � �P ��� � ��  @ �P ��� ���� � �R �P ��� � �@$?   ��j��������� � �P`��� � ���P`��h�� �~�������� � ��P�   ���    �]�����U��S��$�  �ú\  �E�@���E��E�   �E�    �   �E�����    �EЃ��E�E� �E�E����t@���u��u�4���P�ؙ�������u��u�M   �����u䍃h���P貙��������u��u�x���P蘙�����E��E��E�;E��j������]�����U��S��$��  ���[  �E������    �EЃ��E���E� ���E���h�� �<������E� %   ��t���E� ����E���h�� �������E� %   ��uӋE� �E��E�����u���u��u������P�Ę�����0  ���u�u�'  ���E�}� t���u������P萘������   ��jj �E�P�C������E�Pj�u�u�  ���E�}� t���u�����P�F������   �E���%�   �E��E����E�����RP��P���P�������E�����P��x���P����������u荃����P�������}� u)���u������P�Ɨ������������P贗�����#�}�u�������P蚗�����}�	u�  �]�����U��S��$��  ���Y  �z������ � �E�E��@�E���E��E���E��E���E��E�f�@  �E�f�@  �E�E�f�P��� � �E���` � �E���` � �E��� � � �E���u�jjj �u��u��B  �� ��j jjjj�u��*  �� ��j@j j jj �u�j �u��u��  ��0�U��E�P8���u�j��������u���  ���E����u�������E�@8   �E��]�����U��S��$��  ���X  �H������ � �E���` � �E��� ` � �E���` � �E��� � � �E���� � �E���� � �E܋E��@�E�� �Ȁ�E܈�E�f�@  �E�E�f�P�E�f�@ �E���u�Pjj �u��u��	  �� �E���uPjj�u��u���  �� ��j j j jj�u���  �� �E��j@j Pjj �u��u��u��u��X  ��0�U�E�P8���u���������u��  ���E؃��u�'������E�@8   �E؋]�����U��S��4�k  ��kW  �E�E��������� � �E�E��@	�E���E��E���E��E���E��E�f�@  �E�f�@  �UԋE�f�P��` � �E��� � � �E���� � �E���` � �E���u�jjj �u��u��  �� ��j jjjj�u��  �� �E��j@j Pjj �u�j �u��u��  ��0�U�E�P8���u����������u��R  ���E����u��������E�@8   �E��]�����U��S���2  ��2V  ��� � �@$�E�E����t�������P臓������   �E����t?����H���P�f�������� � �P$��� � ��߉P$��� � �@$   �   �E����t����k���P�������l�E����t��������P��������N�E����t��������P�������0�E�� ��t��������P�Ò������������P诒������� � �U�P$��]�����U��S���
  U  �E�'  �U�R�U��U�����t���� ���R���X������   �   �U�����t����P���R���0������   �   �U���@��t��������R���������   �c�U��� ��t��������R���������   �>�U�J��M��u��������R��軑�����    ��U���   ���$����    �]�����U���  T  �U�E��E�@   �} u�E���E��	��  �E�P�H�}u�E���E��	��  �E�P�#�}u�E���E��	��  �E�P�U�E�P�E�@     �]���U����c  _S  �E(���E��	E$��	�E ��@�E��E�   @�} u�M�   P�} t�M��E���E��E�U��P�E�U��P�U�E�P�U�E�P�E�@   �E�@    �E���E��E�U��P�E�@�̀�E�P�E�U��P�E�@    �E�@   �E�@   �E�@@   �����U��WVS��L�i  ��iR  ��������P�֏������j	j �E�P莈������� � �U�Rj	j h )  jh�   jP��  �� �E����E��E����E����E����E����E������u�WVQRP�����P�U����� �E����E�����RP��V���P�3�������� � j j j jj	j jP�C  �� �E�   �9���u䍃r���P���������� � j j �u�jjj#jP�  �� �E��E���9E�~��E�   ��  ��� � j j �u�jjj#jP��  �� ��t
�    �  ��h@B 荄������� � �U�Rj�u�j j h�   jP�  �� �EЃ����;  �EЃ�P�u�������P�0������EЃ����   ��������P��������jj �E�P�Ȇ������� � �U�Rjj h   jh�   j P�  �� �E����E����E����E�����VQRP������P褍���� �E����E����E���QRP�� ���P�}������E����E����E���QRP��4���P�V������E����E����E����E�����VQRP��d���P�$����� �-��������P��������EЃ�P�u�������P��������E��E���9E��'����    �e�[^_]���U��S��$�?  ��?O  �������� � �E�E�E�P�E�E��E�E�f�P�E �E�f�P�E�E�f�P��` � �E��� � � �E���� � �E���` � �E���u�jjj �u��u������� �E ���u$Pjjj�u��~����� �E��j@j Pjj �u�j �u��u�������0�U�E�P8���u���������u��5������E����u��������E�@8   �E��]�����U��S���  ��N  ��� � �E���` � �E���` � �E��y����E��    �E��@   �E�@�U��	E�P�E�@   ��E�P�E�@��E�P�E�@���E�P�E�@���E�P�U�E�P�E��@   �U�E��P�E���E���E��@   �E��@��@�E��P�E��@   �E��P�E��@�� �E��P�E��@���E��P�E��P�E	E��P�E��@   @�E��@   �E��@   �E����E��E��@    �E��@ �  �E��@@   �U�E�P8�E�@ �� �E�P ���u��o������E�E�@ ��߉E�P �E�@8   �E�]�����U��S���L  ��LL  ��` � �E���� � �E���` � �E������E��    �E��@   �E�@�U��	E�P�E�@��E�P�E�P�E�P�E�@���E�P�U�E�P�E��@   �U�E�P�E����E��E��@    �E�@   �E�P�E�@�� �E�P�E�P�E	E�P�E�@���E�P�E��@   @�E��@   �E��@   �E���E���E��@    �E��@ �  �E��@@   �U��E�P8�E�@ �� �E�P ���u���������E�E�@ ��߉E�P �E�@8   �E�]�����U��S��$�
  �ìJ  �E�uPjj j j0�u�u�=����� �E�}� t��������P�������    ��  ���u�L~�����E���uj �u�萀�����u�u��u�u�
������E�}� t�������P薇�����    �d  �E�E�E��@�ЋE� ��RP��0���P�c������E� =USBS��   ��h   �}�����E��u�u�j�u�������E�}� t����T���P�������    ��   �E�E��������P��������E� =USBSt��������P�҆�����    �   �E��@����P������P諆�����E��@��t��������P莆�����    �_�E�@��tR�E�@��P������P�d������E�    �%�U��E��� ����P�����P�:������E��}��  ~����E�]���f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f��$Ë$Ë$Ë$Ë<$�                                                ~ � � � � � � � � ~             ~ � � � � � � � � ~                 l � � � � | 8                   8 | � | 8                   < < � � �   <                < ~ � � ~   <                      < <              � � � � � � � � � � � � � � � �           < f B B f <           � � � � � � � � � � � � � � � �        2 x � � � � x             < f f f f <  ~               ? 3 ? 0 0 0 0 p � �              c  c c c c g � � �               � < � < �             � � � � � � � � � � �               > � >                  < ~    ~ <                f f f f f f f   f f              � � � {                | � ` 8 l � � l 8  � |                       � � � �              < ~    ~ <  ~              < ~                           ~ <                      �                         0 ` � ` 0                         � � � �                       ( l � l (                      8 8 | | � �                   � � | | 8 8                                                 < < <                  f f f $                             l l � l l l � l l           | � � � |   � � |               � �   0 ` � �             8 l l 8 v � � � � v           0 0 0 `                             0 0 0 0 0 0               0         0                   f < � < f                         ~                                    0                     �                                                           0 ` � �             8 l � � � � � � l 8              8 x       ~             | �    0 ` � � �             | �   <    � |               < l � �                 � � � � �    � |             8 ` � � � � � � � |             � �     0 0 0 0             | � � � | � � � � |             | � � � ~     x                                                       0                  0 ` 0                      ~     ~                     ` 0      0 `             | � �                       | � � � � � � � |              8 l � � � � � � �             � f f f | f f f f �             < f � � � � � � f <             � l f f f f f f l �             � f b h x h ` b f �             � f b h x h ` ` ` �             < f � � � � � � f :             � � � � � � � � � �             <         <                   � � � x             � f f l x x l f f �             � ` ` ` ` ` ` b f �             � � � � � � � � � �             � � � � � � � � � �             | � � � � � � � � |             � f f f | ` ` ` ` �             | � � � � � � � � |           � f f f | l f f f �             | � � ` 8   � � |             ~ ~ Z       <             � � � � � � � � � |             � � � � � � � l 8              � � � � � � � � � l             � � l | 8 8 | l � �             f f f f <     <             � � �   0 ` � � �             < 0 0 0 0 0 0 0 0 <               � � � p 8                 <         <          8 l �                                                   �       0                                     x  | � � � v             � ` ` x l f f f f |                   | � � � � � |                < l � � � � v                   | � � � � � |              6 2 0 x 0 0 0 0 x                   v � � � � � |  � x       � ` ` l v f f f f �                 8      <                        f f <       � ` ` f l x x l f �             8         <                   � � � � � � �                   � f f f f f f                   | � � � � � |                   � f f f f f | ` ` �             v � � � � � |                � v f ` ` ` �                   | � ` 8  � |              0 0 � 0 0 0 0 6                    � � � � � � v                   � � � � � l 8                   � � � � � � l                   � l 8 8 8 l �                   � � � � � � ~   �             � �  0 ` � �                 p                                        p         p           v �                                    8 l � � � �                 0  @          ===============================================
 %s
 VBE video mode: %dx%dx%d
 GDT and IDT install
 Reading the kernel.bin
 r kernel.bin error read kernel.bin
 x86_64 hardware not supported
 Enable 4-level paging
   %%  �B���B���B���B���B���B���B���B���B���B���B���A��B���B���B���B���B��B���B���B���B���B���B���B���B���B���B���A���B��@B���B���B���B��Divide error
 Debug exception
 NMI Interrupter
 Breakpoint
 Overflow
 BOUND Ranger exception
   Invalide opcode (Undefined opcode)
 Device not avaliable (Not Math coprocessor
)    Double Fault (Erro de codigo)
  Coprocessor segment overrun (reservado)
    Invalide TSS (Erro de codigo)
  Segment not present (Erro de codigo)
   Stack segment fault (Erro de codigo)
   General protetion (Erro de codigo)
 Page fault (Erro de codigo)
 Intel reserved do not use 15
  x87 FPU Floating-Point error (Math fault)
  Alignment check (Erro de codigo)
 Machine check
    SIND Floating-Point exception
 Virtualization exception
 Intel reserved do not use 21
 Intel reserved do not use 22
 Intel reserved do not use 23
 Intel reserved do not use 24
 Intel reserved do not use 25
 Intel reserved do not use 26
 Intel reserved do not use 27
 Intel reserved do not use 28
 Intel reserved do not use 29
 Intel reserved do not use 30
 Intel reserved do not use 31
  CR2 = 0x%x, CR3 = 0x%x, CR4 = 0x%x
 Unclassified Mass Storage Controller Network Controller Display Controller Multimedia Controller Memory Controller Bridge device    Simple Communication Controller Base System Peripheral Input Device Controller Docking Station Processor Serial Bus Controller Wireless Controller Intelligent I/O Controllers  Satellite Communication Controller Encryption Controller Signal Processing Controller Processing Accelerator Non-Essential Instrumentation Co-Processor Unassigned Class (Vendor specific) Non-VGA-Compatible devices VGA-Compatible Device SCSI bus controller IDE controller (ISA Compatibility mode-only controller) IDE controller (PCI native mode-only controller)    IDE controller (ISA Compatibility mode controller, supports both channels switched to PCI native mode)  IDE controller (PCI native mode controller, supports both channels switched to ISA compatibility mode)  IDE controller (ISA Compatibility mode-only controller, supports bus mastering) IDE controller (PCI native mode-only controller, supports bus mastering )   IDE controller (ISA Compatibility mode controller, supports both channels switched to PCI native mode, supports bus mastering ) IDE controller (PCI native mode controller, supports both channels switched to ISA compatibility mode, supports bus mastering ) Floppy disk controller IPI bus controller RAID bus controller ATA Controller (Single DMA) ATA Controller (Chained DMA)  Serial ATA controller (vendor specific interface)   Serial ATA controller (AHCI 1.0 interface)  Serial ATA controller (Serial Storage Bus) Serial Attached SCSI (SAS)   Serial Attached SCSI (Serial Storage Bus)   Non-Volatile Memory Controlle (NVMHCI)  Non-Volatile Memory Controlle (NVM Express) Other mass storage controller Ethernet controller Token ring controller FDDI controller ATM controller ISDN controller WorldFip Controller PICMG 2.14 Multi Computing Infiniband Controller Fabric Controller Other Network controller  VGA Compatible controller (VGA Controller)  VGA Compatible controller (8514-Compatible Controller ) XGA controller  3D controller (Not VGA-Compatible) Other Display controller Multimedia video controller Multimedia audio controller (AC'97) Computer telephony device   Audio Device (Intel High Definition Audio (HDA) Controller) Other Multimedia controller RAM controller FLASH controller Other Memory controller Host bridge ISA bridge EISA bridge MCA bridge   PCI-to-PCI Bridge (Normal Decode)   PCI-to-PCI Bridge (Subtractive Decode) PCMCIA bridge NuBus bridge CardBus bridge    RACEway bridge (Transparent Mode)   RACEway bridge (Endpoint Mode)  PCI-to-PCI Bridge (Semi-Transparent, Primary bus towards host CPU)  PCI-to-PCI Bridge (Semi-Transparent, Secondary bus towards host CPU) InfiniBand to PCI host bridge Other Bridge Serial controller (8250-Compatible (Generic XT))    Serial controller (16450-Compatible )   Serial controller (16550-Compatible )   Serial controller (16650-Compatible )   Serial controller (16750-Compatible)    Serial controller (16850-Compatible)    Serial controller (16950-Compatible)    Parallel Controller (Standard Parallel Port)    Parallel Controller (Bi-Directional Parallel Port)  Parallel Controller (ECP 1.X Compliant Parallel Port)   Parallel Controller (IEEE 1284 Controller)  Parallel Controller (IEEE 1284 Target Device) Multiport Serial Controller Modem (Generic Modem) Modem (Hayes 16450-Compatible Interface)    Modem (Hayes 16550-Compatible Interface)    Modem (Hayes 16650-Compatible Interface)    Modem (Hayes 16750-Compatible Interface)    GPIB (IEEE 488.1/2) Controller Smart Card   Other Simple Communication controller PIC (Generic 8259-Compatible) PIC (ISA-Compatible) PIC (EISA-Compatible)  PIC (I/O APIC Interrupt Controller) PIC (I/O(x) APIC Interrupt Controller)  DMA controller (Generic 8237-Compatible)    DMA controller (ISA-Compatible) DMA controller (EISA-Compatible)    Timer (Generic 8254-Compatible) Timer (ISA-Compatible) Timer (EISA-Compatible) Timer (HPET) RTC (Generic RTC) RTC (ISA-Compatible) PCI Hot-plug controller SD Host controller IOMMU Other System peripheral controller Keyboard controller Digitizer Pen Mouse controller Scanner controller Gameport controller (Generic)  Gameport controller (Extended) Other input controller Generic Docking Station Other type of docking station 386 486 Pentium Alpha Power PC MIPS Co-processor    FireWire (IEEE 1394) controller (Generic)   FireWire (IEEE 1394) controller (OHCI) ACCESS Bus SSA USB (UHCI Controller) USB1.1 (OHCI Controller) USB2.0 (EHCI Controller) USB3.0 (XHCI Controller) USB Controller (Unspecified )    USB Device (Not a host controller) Fiber Channel SMBus InfiniBand IPMI Interface (SMIC) IPMI Interface (Keyboard Controller Style)  IPMI Interface (Block Transfer) SERCOS Interface (IEC 61491 CANbus iRDA controller Consumer IR controller RF controller Bluetooth Controller Broadband Controller   Ethernet Controller (802.1a – 5 GHz)  Ethernet Controller (802.1b 2.4 GHz)    Other type of wireless controller I2O Satellite TV controller Satellite audio controller Satellite voice controller Satellite data  controller  Network and Computing Encrpytion/Decryption Entertainment Encryption/Decryption Other Encryption/Decryption DPIO module Performance counters Communication synchronizer Signal Processing Management    Other Signal Processing Controller Null PCI Listing devices:
 %s , B%d:D%d:F%d
 Other PCI Device ClassCode (%X), B%d:D%d:F%d
   panic: RAID Controller
 IDE Controller not found!
 RAID Controller not found!
 AHCI Controller not found!
 Uinidade%d PATA
 Uinidade%d PATAPI
 Uinidade%d SATA
 Uinidade%d SATAPI
 Uinidade%d Not found
    e��,c���d��d��e��PANIC,ATA Modo CHS not suport Unidade%d
    Initializing the ATA Controller:
   PIC: Massa Storage Controller not found!
   PANIC: IDE/AHCI PCI Configuration Space
 IDE Controller:
 AHCI Controller:
 IDE or AHCI controller not found    SATA SATAPI SEMB PM sata(x) Read disk CMD ATA IDENTIFY error
 port(x) is hung 
 sata(x) read disk CMD ATA IDENTIFY error
   sata(x) read disk CMD ATA IDENTIFY error ---
 sata%d device not found
 sata%d device type: %s
 Default Unknown IntelliMouse                      1234567890-=	qwertyuiop[]
 asdfghjkl;'` \zxcvbnm,./                                                                                                                                                                                                           !@#$%^&*()_+	QWERTYUIOP{}
 ASDFGHJKL:"~ |ZXCVBNM<>?                                                                                                                                                                                                          [EHCI] Reset of EHCI Host Controller is succeed.
 EHCI initialize
  PCI PANIC: EHCI (USB2.0) Controller not found!
 vid 0x%x, did 0x%x, mmio 0x%x
  Host Controller Initialization
 [EHCI] Port %d : connection detected! Port info %x
 Port info %x
   [EHCI] Port %d : no connection! Port info %x
   [EHCI] Port %d : Port is not enabled but connected, portifo %x
 [EHCI] Port %x : Unable to set device address...
   [EHCI] Port %x : Unable to get devicedescriptor...
 Magic number at descriptor (0x%x 0x%x)
 Max Packet Size %x 
 Device Class %x 
  [ECHI] Port %x : No class found! Asking descriptors...
 Nelson, tem que configurar o dispositivo
 USB Class Mass Storage
   [EHCI] Interrupt: transaction completed
    [EHCI] Interrupt: error interrupt
 [EHCI] Interrupt: portchange
    [EHCI] Interrupt: frame list rollover
  [EHCI] Interrupt: host system error
    [EHCI] Interrupt: interrupt on advance
 [EHCI] Interrupt: unknown
  [EHCI] Transmission failed due babble error
    [EHCI] Transmission failed due transaction error
   [EHCI] Transmission failed due serious error
   [EHCI] Transmission failed due data buffer error
 EHCI FAIL Timeout
    USB HUB install
    Hub descriptor: len:%d, typ:0x%x, cnt:%d, char:0x%x, pwg:%d, curr:%d
 hubdesc.variable[] = %x,%x
 Power on - port %d
   Hub Port%d A device is present on this port, status: %x
 PORT_ENABLE
   length %x, type 0x%x, bcdusb 0x%x, class 0x%x
  subclass 0x%x, protocol 0x%x, maxpacketsize 0x%x
   vendorid 0x%x, productid 0x%x, devicever 0x%x
  vendorstr 0x%x, productstr 0x%x, serialstr 0x%x,   				confcount 0x%x
 PORT_DISABLE
    Hub Port%d No device is present on this port, status: %x
 [SMSD] Sending bulk error
 [SMSD] Recieving bulk error
   csw->signature %x, csw->status %x
  [SMSD] Recieving command status wrapper error
 [SMSD] Status at end
    [SMSD] Command Status Wrapper has a invalid signature
 [SMSD] Status=%x 
 [SMSD] Status is not 0 
 [SMSD] Data residu %x 
 %x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �� �� �� ̱ ر � ��  � P� p� �� �� � � 0� M� l� �� �� ̳ � � #� A� _� }� �� �� ״ �� � 1� t� �� �� �� �� յ � �� � /� G� W� a� w� �� �� ˶ � �� �                                                                                                                                                                                 3�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         @�     c�    ~�    ��   ��  � 
 �  |� � � � 4� � �� �  �   ��   ��   ��   �� 0 ں   ��  ,�  X�   ��  ��  ̻  ��  �  �    >�   R�   h�   x�   ��   ��   ��   Ƽ   ܼ  � �    �   4�   l�   |�  � ��    ��   Խ   ��   �  � P�    l�   {�  � ��    ��   ��   ��   Ǿ   Ծ  ��   �   -�   :�   L�  p� @	 �� �	 Կ  
 �  � 7�    D�   x�   ��   ��   ��   �   @�   h�  ��  ��  � � 0�   ^�   z�  ��  ��  ��  �   @�   _�  � l�    ��   ��   ��   ��     �   (�  T�  t�   ��  ��  ��  ��   ��  �   �   3�   F�  � L�   	 o�  	 ��  	 ��  	 ��  	 �� 	 ��  �	 ��   
 
�  �
 "�    @�   D�   H�   P�    V�  0 _�  @ d�    t�   ��   ��   ��   ��  ��   � 0 � � 7� � X�   {�   ��   ��   ��  ��  ��   ��  	 �    �   /�   F�   T�   i�    ��  ! ��  � ��    ��    ��   �   )�   D�    `�   ��  � ��    ��   ��   ��    �  � (�     K�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     t� y� �� �� O� W� W� _�                     S1 �{ S1 S1 S1 S1 S1 S1 S1 S1 S1 g1 �w S1 S1 S1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        zR |�  4      �����   H Gu Duxu|�� A�A�C      T   ���          h   '���A    E�By�     �   x��          �   4���    E�BW�     �   3���3    E�Bk�     �   F���    E�BL�      �   :���   E�BD����       ���   E�B�   @  	���F    E�B~�     `  /���Q    E�BI�    �  `���T    E�BL�    �  ����2    E�Bj�      �  �����   E�BD����   �  x���A    E�By�       ����g    E�B_�     $  ����m    E�BD�a��     H  )���}    E�BD�q��    l  �����    E�B�� ,   �  ���\   E�BF���K�A�A�A�       �  8���*    E�BD�^��      �  >���`    E�BD�T��       z���n    E�BG�_��     (  Ċ��D    E�BD�x��      L  ���*    E�BD�^��     p  ���K    E�BC�    �  ����    E�B��    �  ����&    E�B^�      �  �����    E�BD����    �  n����    E�B��      ���          (  Č��H    E�B@�     H  ����   E�BG����,   l  �����   E�BF���o�A�A�A�       �  ����    E�BD����     �  �����    E�BD���� ,   �  r���g   E�BF���V�A�A�A�         ����s    E�BD�g��    8  ����E    E�B}�     X  ���E    E�B}�      x  L����   E�BD����   �  ���^    E�BD�    �  &���q   E�BD�e��   �  s���    E�BL�      �  g���#    E�BD�V�A�       f���U    E�BM�    @  ����~    E�Bv�    `  ����|    E�Bt�    �  U���`    E�BX�    �  ����Y    E�BQ�    �  Μ��`    E�BX�    �  ���Y    E�BQ�        G���=   E�BD�1��   $  `����    E�B��    D  ����    E�B��    d  Ο���    E�B��    �  �����    E�B��    �  e���"    E�BZ�     �  g���"    E�BZ�     �  i���*    E�Bb�       s����    E�B��    $  ���:    E�Br�     D  ���G    E�B�     d  (���G    E�B�     �  O���E    E�B}�     �  t���E    E�B}�      �  ����J    E�BA�A��     �  ����{    E�BD�n�A�    	  ���:    E�BA�p�A�     0	  ,���:    E�BA�p�A�     T	  B����   E�BD����    x	  ����    E�BA���A�    �	  h����   E�BD����    �	  /���c   E�BD�W��    �	  n����   E�BD����    
  ���j   E�BD�^��    ,
  K����   E�BD����    P
  ݱ��N   E�BD�B��    t
  ���m    E�BD�a��    �
  P���W    E�BO�    �
  ����F    E�B~�      �
  �����    E�BD���� ,   �
  7���}   E�BF���l�A�A�A�      ,  �����    E�B�� ,   L  ���_   E�BF���N�A�A�A�   ,   |  ���   E�BF�����A�A�A�       �  ���;   E�BD�/��   �  
����    E�B�� ,   �  r���S   E�BF���B�A�A�A�   ,      ����d   E�BF���S�A�A�A�   ,   P  ����D   E�BF���3�A�A�A�   ,   �  ����D   E�BF���3�A�A�A�      �  X��       (   �  �����    E�BF�����A�A�A�(   �  �����    E�BF�����A�A�A�     K����    E�B��     <  ����@    E�BD�t��  $   `  ����   E�BE����A�A�(   �  �����   E�BE��}�A�A�       �  -���   E�BD����     �  ����    E�BD���� (   �  �����    E�BF�����A�A�A�(   (  ���Q    E�BF���@�A�A�A�(   T  B����    E�BF�����A�A�A�$   �  ����)    E�BB��]�A�A� (   �  ����T    E�BF���C�A�A�A�   �  ���+    E�Bc�     �  ���M    E�BE�       E���0    E�BD�d��     8  Q���    E�BR�     X  K���    E�BU�     x  H���    E�BW�  ,   �  G����   E�BF�����A�A�A�      �  D ��           �  �����    E�BD����       ����    E�Bz�       ����z    E�Br�    @  ;���'    E�B_�      `  B���Q    E�BD�E��     �  o���8    E�BD�l��     �  ����J    E�BB�     �  ����z   E�BD�n��$   �  ����   E�BD���A�   $     ����-   E�BA�#�A�       <  ����8    E�BD�l��      `  ����:    E�BD�n��     �  ����J    E�BB�     �  ����*    E�BD�^��      �  �����    E�BD���A�    �  �����    E�BD����      U���F    E�B~�     0  {���5    E�Bm�     P  ����5    E�Bm�     p  ����%    E�B]�     �  ����%    E�B]�     �  ����4    E�Bl�     �  ����%    E�B]�      �  ����v    E�BD�j��       ����    E�BD����     8  ����s   E�BD�g��    \  �����    E�BD����     �  �����   E�BD����    �  S���2   E�BD�&��    �  a���X   E�BD�L��    �  ����9   E�BD�-��      ����,   E�BD� ��    4  ����   E�BD����    X  �����    E�B��    x  ����    E�B�� ,   �  ����,   E�BF����A�A�A�       �  ����*   E�BD���    �  �����   E�BD����      �����   E�BD����    4  ���   E�BD���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            GCC: (Ubuntu 9.3.0-17ubuntu1~20.04) 9.3.0                                    �           �           �           �           �            �            �            �      	     ��      
      �            �                                 ���             8           �        $    p        +            ��2            ��9            ��B            ��K            ��Q            ��\            ��d            ��o   �  H     y   �"        }   �"        �   �!        �   "        �   �!        �   @"        �            ���   $# �    �            ���   Z' g    �            ���   �)        �   �+        �            ���            ���   �� @    
 �            ��3            ���   �< �      i@ �     %  A �    4  �B c    H  VE �    b  E        g  ,C        l  �D        q  D        v  E        {           ���  �Z �     �  �O W     �  CP F     �  �P �     �  7Q }    �  �S �     �  @T _    �  �U     �  �W ;    
  f[ S      �] d               ��)           ��.           ��6           ��<           ��E           ��Q           ��W           ��]           ��e  0�      u  4�      �  p      �  �y -    �           ���  p      �  p      �           ���  2 �     �           ���           ��             ���   �          �        � *       >*       $  ۑ �    6  � T     =  u z     G  8 �     _  � n     ]  8! �    f  �{ *     w  `< :     �  �x      �  A,       �  ��      �  ��      �  �; {     �  e+       �  �*       �  �      �  hl )     �  K4 =    �  �w �      �,       
  � �       >~ %     5  p      =  +       C   �      G  �*       M  ��      X  n,       ^  ��     	 h  �,       n  {9 �     w  �( s     �  ��      �  *       �  �1 ~     �  _,       �  �j �     �  �      �  �% �     �  6� �     �  { :     �  � Q     �  P,         )+         y) E       �+         (�      !  �+       '  ,�      /  S1      ;  g1 #     I  " `     N  /9 "     _  ; E     l  �u Q     x  <p      �	  � 3       ��  @    �  p      3
  {J �    �  z       �   � �    	 �  �+       �  �5 �     �  �      �  �      �   p      �  $p      �  A        �        +       
  u }       ]m 0     =  �      A  },       G  Hp 
     M  t+       S  /*       Y  /v J     h  �3 `     ~  Tp      �   �       �  �t �     �  �� �     �  �| �     �  �} 5     �  � g     �  �      �  �      �  ,       �  �*       �  ~ %       �: G     %  �� �    4  �� 9    R  �{ �     c  I: G     u  �*       {  : :     �  X6 �     �  93 Y     �  �x      �  �s �     �  �1 U     �  �� 2    �   *       �  � �       �2 `       (p      x  ]       #  Te     �   �       8  *       >  ��      I  ��     	 Y  � �     �  Dp      r  � A     _   �      h  &< :     �
   �       u  �x      �          �   �       G
  �z      �  �m      �  �k �     �  �� *    �   �  �    7
  �c �     �  � �     �  lp 
     �  V+       �  ` A     �  �*       �  �u 8     	  Yf �    �
   �       	  � \    	  �/ q    %	  ,       +	  �, �    >	   �      �
  I j    T	  ,p      ]	  0p      f	   `      j	  �i �     u	  �m �    �	  �x      �	  ]2 |     �	  f  �     �	  �m      �	  �h     �	  �,       �	  �*       �	  �/ ^     �	  � D     F
   �       �  M F     �	  u '     �	  � �    �	  xp      �	  i} F     �	  ��      �	  Q &     �   p      
  ��     	 
  a; J     
  �� ,    +
  4 *     2
  aa D    D
   �       K
  Ik Q     X
  4) E     ]
  8+       c
  �*       i
  �l +     p
  �z 8     �   �p      ~
   �      �
  k*       �  p      �
  �~ v     �
  yv z    �
   �       �
  �+       �
  w �     �
  $�      �
  �} 5     �
  D�     �
  ` D    �
  `        �x 
       p      $  \*       *  8�      E
   �       0   m     �  ��      =  `      A  �~ %     d  Q9 *     m  m M     t  �m      �  �*       �  :     �  O m     �  67 �     �  -� X    �   �       �  �)       �  1L N    �  ^ K     �  j �    �  '       �          �  M*         �*       	  @p        `        ��        9 "     ,  �+       2   p      @  8,       F  �� ,    S   �      X  �*       ^  �x      l  & �     �  �*       �  ),       �  � s    �  u*       �  O       �  �+       �  c~ 4     �  8 2     �          �  kd �     �          �  4p      �  8p      �  e @       ��     	   �,       %  �l T     2  G+       8  �x      C  ��      T  �     m  �      r  ;{ J     �  �3 Y     �  �: E     �
  �b �     �  &       stage2.asm gdt_flush.flush start64 _stack main.c data.c stdlib.c string.c gui.c font8x16.c stdio.c vsprintf.c _vsputs_r .L8 .L9 .L14 .L13 .L12 .L11 gdt.c set_gdt idt.c set_gate_idt vetor.asm isr_jmp irq_jmp exception.c irq.c fnvetors_handler pci.c ata_pci_configuration_space ata_bus_install detect_devtype ata_identify_device set_ata_device_and_sector .L57 .L56 .L55 .L54 .L52 ahci.c sata_port_initialize stop_cmd start_cmd sata_port_confg sata_set_cfis sata_set_prdt sata_set_cmdHeader ahci_ata_indentify sata_identify ahci_read ahci_write storage.c fs.c cpuid.c msr.c paging.c bootblock.c pic.c ps2.c mouse.c largura_da_tela altura_da_tela status.1173 mouse_refresh keyboard.c shift caps_lock ehci.c ehci_pci_configuration_space bulk.c hub.c _GLOBAL_OFFSET_TABLE_ __x86.get_pc_thunk.cx putchar isr05 ehci_recieve_bulk strcpy kbdc_wait pci_scan_bcc_scc_prog vsprintf keyboard_install ata_pio_write ata_record_channel irq07 mouse_x count_mouse ata_soft_reset isr27 isr13 __x86.get_pc_thunk.di cpuid pci_get_info mouse_handler irq12 ehci_int_td ehci_periodic_schedule_disable ata_pci isr22 td2 isr15 key_buffer irq10 ahci_type irq14 ata_wait idt_install ascii_minusculas isr02 irq_enable irq09 file_read_block initialize_heap gdt_install ehci_sondagem keyboard_write memcpy irq08 isr23 interrupter irq02 pae_pde isr29 pae_pte default_irq irq11_handler puts pci_check_vendor ata_wait_drq mouse_write dv_uid fs_directory mouse_position file_sector_count exception_mensagem isr31 pci_scan_bcc __x86.get_pc_thunk.ax ATA_BAR1 ATA_BAR4 itoa qh1 isr21 clears_creen load_pae_page_directory_pointer_table td3 irq11 gdtr1 isr28 isr04 MOUSE_BAT_TEST pci_read_config_dword gdt2 eh_frame pic_install ehci_init_qh ehci_memset ehci_start put_pixel_buff ehci_driver __x86.get_pc_thunk.dx irq04 isr20 ehci_periodic_schedule_enable ata_wait_busy ehci_send_bulk ehci_set_device_configuration keyboard_handler ata_wait_not_busy isr14 ata_status_read pci_scan_class write_pci_config_addr dmaphys cof_bootblock irq_function ehci_set_device_address isr03 ehci_port_init read_pci_config_addr CPUID_REQUEST read_directory_entry isr01 first_time pci_class_names fseek font8x16 ata_pio_read ata_record_dev __end load_pml4_table cpuid_processor_brand usb_control_msg ehci_pool draw_char_transparent gdtr2 isr26 put_pixel isr11 mouse_read open_file_r glyph irq_install irq03 exceptions_install __x86.get_pc_thunk.bx ATA_BAR0 ATA_BAR3 qh3 file_close page_install HBA_BASE irq_disable fread enable_pae open_file irq13 isr12 fault_exception fopen kbdc_set_cmd main gdt1 ehc_malloc buttons ftell pci_classes ata_cmd_write usb_hub_init fclose sata_write_sector __data cpuid_vendor trap isr24 isr16 getmsr keyboard_read pml4e isr08 ehci_reset mouse_install __bss irq01 fgetc pdpte ehci_stop usb_stick_send_and_recieve_scsi_command sata_read_sector ehci_pool_start idtr keyboard_charset isr07 speed refresh_rate td1 ehci_asynchronous_schedule_disable pci_size setmsr page_enable isr18 i2hex ahci_initialize pci_scan_bcc_scc ehci_get_device_descriptor isr00 ata_initialize rewind initialize_gui gdt_flush isr06 isr10 dv_num qh2 mouse_y pci_scan_vendor irq00 periodic_list irq06 ehci_handler ehci isr17 hba_mem_space gdt_execute_long_mode isr19 irq05 ehci_init isr09 idt_flush isr30 ehci_asynchronous_schedule_enable strlen __code filename_cmp ATA_BAR2 ATA_BAR5 read_super_block id_mouse_strings irq15 cpuid_string isr25 sata_idtfy ascii_maiusculas ehci_wait_for_completion cmd1 KEYBOARD_BAT_TEST pci_write_config_dword ata_wait_no_drq free  .symtab .strtab .shstrtab .text .text.__x86.get_pc_thunk.bx .text.__x86.get_pc_thunk.ax .text.__x86.get_pc_thunk.cx .text.__x86.get_pc_thunk.dx .text.__x86.get_pc_thunk.di .data .got.plt .data.rel.local .data.rel .bss .eh_frame .comment                                                          �                 !          �  �                    =         � �                    Y         � �                    u         � �                    �         � �                    �          �  �  �?                  �          �  �                   �          �  �  �                  �         �� ��  @                   �          �  �   �                �          �  �                     �      0         *                               , �     Z         	              & �                               �3 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ELF          >     @     @       `�         @ 8  @                 @      @      �      �                   �      �A      �A     �k      �                         @E      @E      0       0             Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �    H�  @    H�  0    H�% �A H����    H�%�A H1����   ������H����  �2�����0��  �2�  0�H���H��H��H��H��L��M������SH��H1�H��H�       H��H��H�H�H��   H��   ��[�� �f "�� �f%��"��������UH��AWSH��   ��H�����I���     L�H��H���H��     �   H��     � H��     �    �(   �    H��������H�H��I��H��������H���H���������H�H�     H���������H��     H� �������H�H�     H��H����H�@�������H��H��H���H��� ��H���������H��H��H���H��I��H�fd������H���H��������H�<I�߸    H�u�������H���H� �������H�<I�߸    H�u�������H���H�2�������H�<I�߸    H�u�������H���I�߸    H��)������H���I��H�E/������H���H�D�������H�<I�߸    H�u�������H���H��H���H��I��H�wQ������H���H�X�������H�<I�߸    H�u�������H���I�߸    H�R������H���H��H���H��I��H�X������H���H��H���H��I��H�^Z������H���I�߸    H���������H���I�߸    H�5�������H���I�߸    H�u������H���I�߸    H�b~������H���H�h�������H�<I�߸    H�u�������H���I�߸    H�pH������H���H�y�������H�<I�߸    H�u�������H��ҿ   I��H��������H���H���������H�<I�߸    H�u�������H���I�߸    H�4?������H���I�߸    H�-x������H��ҿ   I��H�_z������H��п   I��H�_z������H��п   I��H�_z������H���H���������H�<I�߸    H�u�������H���I�߸    H��������H���H��`�����   �    H��I��H��������H���H��`���H��I��H�g������H���H��`���H��H���������H�<I�߸    H�u�������H���H���������H�4�    I��H���������H���H�(�������H�H�H�(�������H�H�H���������H�H�H���������H�4�    I��H���������H���H���������H�H�H���������H�H�H���������H�H�H���������H�4�    I��H���������H���H��������H�H�H��������H�H�H���������H�H�H���������H�<I�߸    H�u�������H���H��������H�<I�߸    H�u�������H���I�߸    H���������H���H�*�������H�<I�߸    H�u�������H���I�߸    H���������H���H�6�������H�<I�߸    H�u�������H���I�߸    H��6������H��ҿ   I��H�R�������H���H��     H�H�@�������H�H�H��     H�H�H���������H�H�H��     H�H�P�H�A�������H�<I�߸    H�u�������H���I�߸    H��������H���H��     �H��X���H�¾   �   I��H��^������H���H��������H�H� H��H��X���H�  j j A�    A��   �    H��H�H�������H�H��I��H�Ă������H���H��I�߸    H��N������H��Ҹ    ����H��     ���u��H�G�������H�<I�߸    H�u�������H��ҿ   I��H�R�������H���H�      H�H�      H�H�W�������H�4H��I��H��������H���H�Z�������H�4H�^�������H�<I��H���������H���H�E�H�}� tOH�      H�H�U�H��H�¾    �    I��H���������H���H�E�H��I��H�Ô������H����%H�k�������H�<I�߸    H�u�������H��Ҹ    ��H��     ��PH��     �H��H���H��I��H��B������H��АH�e�[A_]���UH��H����H�����I�n�     L؉}�E�E��怋E��P��U���u�����UH��H��8��H�����I�,�     L�H�}��u�U��M�E��E��D�E�}�u �M(�U0�E8E��D�M�E��D�M�D�E�@�}�@�u؈MԈUЈE̋E�H�H��    H�E�HЋU�������� 	�f�����P�� 	ʈP�E�H�H��    H�E�HЋU������H�� 	�Hf�����P�� 	ʈP�E������E�H�H��    H�E�HЉʈP�E�H�H��    H�E�H��U���у��P���	ʈP�E�H�H��    H�E�H��U���������P���	ʈP�E�H�H��    H�E�H��U����������P��	ʈP�E�H�H��    H�E�H��U܃������P��	ʈP�E������E�H�H��    H�E�Hȃ������B���	ȈB�E�H�H��    H�E�H��U؃��������P���	ʈP�E�H�H��    H�E�H��Uԃ��������P���	ʈP�E�H�H��    H�E�H��UЃ��������P��	ʈP�E�H�H��    H�E�H��Ũ������P��	ʈP�E������E�H�H��    H�E�HЉʈP�����UH��AWS��H�����I�d�     Lۺ   �    H�H     H�<I��H��������H���j j j j j j A�    A�    �    �    �    H�H     H�<H��&������H���H��0j j jj jj A�   A�
   �    �    �   H�H     H�<H��&������H���H��0j j jj jj A�   A�   �    �    �   H�H     H�<H��&������H���H��0j j jj jjA�   A�
   �    �    �   H�H     H�<H��&������H���H��0j j jj jjA�   A�   �    �    �   H�H     H�<H��&������H���H��0H���������H�jj j j jjA�    A�	   ���g   �   H�H     H�<H��&������H���H��0H���������H�H��0��H���������H�H�� j j j j j j A�    A�    �щ¾   H�H     H�<H��&������H���H��0H�(     f�� H�H     H�H�(     H�DH�(     H�<I��H��������H���I�߸    H��,������H��ҿ+   I��H��,������H��АH�e�[A_]���UH��H����H�����I�g�     L؉}��E�f�� ؐ����UH��AWS��H�����I�5�     Lۺh   �    H�H     H�<I��H��������H���H�P�������H�H� H�H     H�D�[A_]���UH��H�� ��H�����I���     L؉}�H�u�D��D��f�U��ʈU���U��U�H�U���H��     �U�Hc�H�H��H��
�� 	�f�
H��     �U�Hc�H�H��H��J�� fM�f�J�U��H��     �M�Hc�H�H��H�փ��Q���	�QH��     �U�Hc�H�H��H��J���J�U�у�H��     �U�Hc�H�H��H�΃��J���	�J�U�у�H��     �U�Hc�H�H��H�������J��	�J�U�у�H��     �U�Hc�H�H��H�����J��	�JH�U�H����H��     �U�Hc�H�H��H��J�� 	�f�JH�U�H�� ��H��     �U�Hc�H�H��HʋJ�� 	�JH��     �U�Hc�H�H��HЋP�� �P�����UH��AWS��H�����I���     Lۺ   �    H��     H�<I��H��������H���I��H�A:������H���I�߸    H��k������H���I��H�Go������H���I�߸    H�?�������H���H��+     f��H��     H�H��+     H�DH��+     H�<I��H��������H��А[A_]���UH��H����H�����I���     L؉}��u�f�U�ʈU��M��U�u��}�j A�   A�ȹ�   I�3-������J���H�������UH��H����H�����I�U�     L؉}��u�D�E�f�U�ʈU�D�E��U�u��}��M�QA�   ��   I�3-������J���H�����f.�      ��AWAVAUATASARAQAPWVUTSRQP�%�A H��$�   �A  �%�A XYZ[\]^_AXAYAZA[A\A]A^A_��H��   H�h    h    ����h    h   ����h    h   �u���h    h   �f���h    h   �W���h    h   �H���h    h   �9���h    h   �*���h   � ���h    h	   ����h
   ����h   �����h   �����h   �����h   �����h    h   �����h    h   �����h   ����h    h   ����h    h   ����h    h   ����h    h   �{���h    h   �l���h    h   �]���h    h   �N���h    h   �?���h    h   �0���h    h   �!���h    h   ����h    h   ����h    h   �����h    h   �������AWAVAUATASARAQAPWVUTSRQPH��$�   ��5  XYZ[\]^_AXAYAZA[A\A]A^A_��H��   H���AWAVAUATASARAQAPWVUTSRQPH��$�   �5  XYZ[\]^_AXAYAZA[A\A]A^A_��H��   Hπ<%hE  ��  �%hE  �% #E �%�"E �%p"E �%�"E �%�"E H�%8"E H�%#E H�%("E H�%h"E H�<% #E H�4%X"E H�,%�"E L�%�"E L�%`"E L�%�"E L�%�"E L�$%0"E L�,%�"E L�4%#E L�<%�"E H1�H��f�%@"E H��f�%(#E H��f�%�"E H��f�%�"E  �H�%�"E H��A     �k����V  H�%�"E "�H�       ���H��A     �C���H1�f�%@"E f��f�%(#E f��f�%�"E f��f�%�"E f��H�,%�"E H�<% #E H�4%X"E H�%8"E H�%#E H�%("E H�%h"E L�%�"E L�%`"E L�%�"E L�%�"E L�$%0"E L�,%�"E L�4%#E L�<%�"E �4%�"E �4%�"E �4%p"E �4%�"E �4% #E �%hE h    h    �]���h    h!   �N���h    h"   �?���h    h#   �0���h    h$   �!��� �<%�)@ ��  �<%hE  ��  �%�)@ �%hE  �% #E �%�"E �%p"E �%�"E �%�"E H�%8"E H�%#E H�%("E H�%h"E H�<% #E H�4%X"E H�,%�"E L�%�"E L�%`"E L�%�"E L�%�"E L�$%0"E L�,%�"E L�4%#E L�<%�"E H1�H��f�%@"E H��f�%(#E H��f�%�"E H��f�%�"E  �H�%�"E ��\  H�%�"E "�H�       ���H1�f�%@"E f��f�%(#E f��f�%�"E f��f�%�"E f��H�,%�"E H�<% #E H�4%X"E H�%8"E H�%#E H�%("E H�%h"E L�%�"E L�%`"E L�%�"E L�%�"E L�$%0"E L�,%�"E L�4%#E L�<%�"E �4%�"E �4%�"E �4%p"E �4%�"E �4% #E �%hE h    h%   �!���h    h&   ����h    h'   ����h    h(   �����h    h)   �����h    h*   �����h    h+   �����h    h,   ������AWAVAUATASARAQAPWVUTSRQP�%�A H��$�   ��5  �%�A XYZ[\]^_AXAYAZA[A\A]A^A_��H��   H�h    h@   ����h    hA   ����h    hB   �u���h    hC   �f���h    hD   �W���h    hE   �H���h    hF   �9���h    hG   �*���h    hH   ����h    hI   ����h    hJ   �����h    hK   �����h    hL   �����h    hM   �����h    hN   �����h    hO   ����h    hP   ����h    hQ   ����h    hR   ����h    hS   �v���h    hT   �g���h    hU   �X���h    hV   �I���h    hW   �:�����UH��AWS��H�����I���     L�H�p�������H��    �   �ƿ    I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H�h�������H��    �   �ƿ   I��H�70������H���H�x�������H��    �   �ƿ   I��H�70������H���H�0�������H��    �   �ƿ   I��H�70������H���H� �������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ	   I��H�70������H���H���������H��    �   �ƿ
   I��H�70������H���H�p�������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H�`�������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ$   I��H�70������H���H�x�������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H�(�������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H�h�������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H�8�������H��    �   �ƿ   I��H�70������H���H���������H��    �   �ƿ   I��H�70������H���H�h�������H��    �   �ƿ   I��H�70������H��А[A_]���UH��AWSH��0��H�����I�g�     Lۉ}̐H���������H�� ��u�H���������H�� �PH���������H��H�(       �E�H�H�H��H��I��H��������H��Ѓ}���    �H�E� �H�E� �H�E�H�E�H��I��H��d������H���H�E�H�E�H�� H��H�M�H�U�H�E�I��H��H��H�P�������H�<I�߸    I�u�������I�A��H�E�H�� H��H�E�H��H��H�y�������H�<I�߸    H�u�������H���H���������H�H� H���   H��H���������H�<I�߸    H�u�������H�������UH��AWH��(��H�����I�ݽ     L�H�}�H�u�H�@�������H�H�H�U�� H�U�H��   H9U�tH�U�H��`  H�U�H�}� u���H�}� tZH�U�H���   H���������H�H�
H�U�H��  H�X�������H�H�
H�U�H��  H��I��H��n������H�����H��(A_]���UH��AWSH��p��H�����I��     L�H�}��E�    H�E�    H�E�    f�E��(   �    H�(,     H�<I��H��������H���H�(,     H�H����  H��    H�)� H�H�� H�>��H�(,     H�DH�E�H�(,     H�D H�E�H�(,     H�D(H�E�H�(,     H�DH�E��H�E�H���������H�4H��I��H���������H���H�E�H�}� uuH�E�H��H���������H�<I�߸    H�u�������H���H�E�H��I��H���������H���H�E�H�E�H��  H�E�H��H��I��H�)�������H����  �E�    H�E�    H�}� tTH�E�� �E�H�E�H�E�H�E�H�E�   �E�    �'�E�H�H��    H�E�H�H�E�H�H�E�   �E��}�~�H�E�H��I��H���������H���H��H�M�H�U�H�uЋE�I����I��H��������H���H��uDH�E�H��I��H���������H���H�E�H�E�H��  H�E�H��H��I��H�)�������H���H�E�H��I��H�Ô������H����E�    �(   �    H�(,     H�<I��H��������H��и    ���  H�(,     H�DH�E�H�(,     H�DH�,     H�H�(,     H�D(H�E��H�E�H���������H�4H��I��H���������H���H�E�H�}� u.H�E�H��H���������H�<I�߸    H�u�������H����UH�U�H�E�H��H�¾    �    I��H���������H���H�,     H�    H�E�H��I��H�Ô������H����E�    �(   �    H�(,     H�<I��H��������H��и    ���H  I�߸    H�K�������H����E�    �%  I�߸    H���������H����E�    �  �H�(,     H�TH�(,     H�D H��H��H�B������H����E�    �(   �    H�(,     H�<I��H��������H��и    ���   �H�(,     H�D H�E�H�E�H��I��H���������H���H�E�H�E�H�ƿ    I��H���������H��к(   �    H�(,     H�<I��H��������H��и    ���E�    ��E���}� u��    �怃E���������UH��AWATSH��X��L�%����I��     M�H�E��  H�E��  �E�    H���������I�<M��    H�u�������L���H� �������I�H�H���������I�H� H��������I�H��H��M��H�	�������L���H�E�H�}� u*H�"�������I�<M��    H�u�������L����g  H�E�H�E�H�E��@��H�E�H�H�E�H�E��@$��H�h,     I��  H�E�,�   H�E�� ����tn����   ��t��t<�wH�E�H��� ������ta�E܍P�U�H�U��RH�h,     H�L��<H�E�H��� ��H�h,     I��	  �H�E�H�@H�h,     I��  ��H�E�H��� ��HE�H�E�H;E��F����E܉�H�h,     A��   �   �����H�h,     A��  H�h,     I��  H�h,     I��	  H�h,     A��   ����H�8�������I�<M��    I�u�������M�A���E�    �DH�h,     �E�H�L������H�k�������I�<M��    H�u�������L��҃E�H�h,     A��   ��9E�|�H�h,     A��  ����H�o�������I�<M��    H�u�������L���H�{�������I�<M��    H�u�������L��Һ   �   � �  M��H�o�������L���H�x�������I�H� H�E�H�E��     H�E��     H���������I�H� H�E��E�    �T  H�h,     �E�H�L��H�h,     A��  8��  ��  H�E��� �  H�x�������I�H��(�  H� �������I�H�H��������I�H� �0�  H��8�  H��N������I�H�H�m�   H�E�H�  �     H�E�H  � %��� �E�����H�E�H  H����	��H�E�H   � %  ����H�E�H   H���Ѐ�ŉ�H�E�H   � %   ��u�H�E�H  � %��� �E�����H�E�H  H����	��H�E�H   � %  ����H�E�H   H���Ѐ̅��H�E�H   � %   ��u�
   M��H��O������L����E�    �   H�E�H�  �     H�E�H  � %��� �E�����H�E�H  H����	��H�E�H   � % �����H�E�H   H����  ���   M��H�P������L����H�E�H   � %   ��u�E��}��]������E�H�h,     A��   ��9E������H�E�� ��H���������I�<M��    H�u�������L���H��X[A\A_]���UH��H����H�����I�0�     L�H�E��  H�E��    �����UH��AWATSH��(��L�%����I��     M܉}��E�    �   ����؉E܃}���   �}��}�t�}��q��  M��H��O������L���H���������I�H� H   �H���������I�H� H�� � ��H���������I�<M��    H�u�������L�������_�����UH��H����H�����I�#�     L؉}��E�    ���E��E�i�'  9E�|퐐����UH��H����H�����I�ܯ     L؉}��E�    ���E��E�i�'  9E�|퐐����UH��H����H�����I���     L� �H�U�H�U�H��H��P������H����E��   ���m��}� �������UH��H����H�����I�;�     L�H�}�H�E�"ؐ����UH��H����H�����I�	�     L�H�}�H�E�"ؐ����UH����H�����I�ۮ     L� ��� "��]���UH����H�����I���     L� �   �"��]���UH��H����H�����I�}�     L�H�}�H�U�H�� ���H�u�H�U�H�h     H�H�U�H��   H��H�p     H�H�U�H��    H��H�x     H�H�U�H�� 0  H��H��     H������UH��AWSH����H�����I�٭     L�H��-     H�   H��-     H��   �    H��I��H��������H���H��-     H�H�E�H��������H�H� H������H��������H�H� H������H��������H�H� H������H�E�H��H��H��������H�H� H��H������   H!�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH��-     H�    �H��[A_]���UH��AWSH��`��H�����I�:�     L�H�}�H�u��U��M�H��-     H�H�E�H��-     H�HA  H��H�E�H�E�H�E�H�E�H�E�H��-     H��E��}�   @v:H���������H�<I�߸    H�u�������H���H�E�H�     �   �  �   +E���9E�vN�   +E������E���H���������H�<I�߸    H�u�������H���H�E�H�     �   �-  �E����E܋E�%�  ��t�E��E܍��  ��H���	�E؋E�%�  ��t�E��E�H�����H�E��    H��I��H��������H����E�    ��   H�E�����H�E�����H�E������E�����tH�E�����H�E�H��H��H������   H!�H�E�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH�E�H�E�   �E��E�;E�����H�E�H�E��E�    �r  �U��E��H�H��    H�E�H������U��E��H�H��    H�E�H������E�����t!�U��E��H�H��    H�E�H������U��E��H�H��    H�E�H�����H�E�H��H���U��E��H�H��    H�E�H�H������   H!�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH�E�   H��-     H�H�PH��-     H��E��E�;E������I�߸    H�_P������H��ҋE���-   @��H�E�H��    H��`[A_]���UH��AWSH�� ��H�����I�ߧ     L�H�}�H��-     H�   �E�   �U�H��-     H������H��I��H��������H��ЋE�E��E� 8  �E�H��-     H��U�Hc�Hщ¾    H��I��H��������H���H��-     H�H�� [A_]���UH��AWH��(��H�����I��     L�H��-     H�H   H�E��E� � �E��  �r�E�    �ZH�E�� ���E�����������u<H�E�� �ƋE�   �����	���H�E��E��    �E�� @  �����C�E��}�~�H�E��E��E�9E�r�H��������H�<I�׸    H�u�������H������H��(A_]���UH��H��(��H�����I�!�     L�H�}�H�U�H���U��U����U��U����U�H��-     H��E�H�H�E�H�E�� �E��   �������!Љ�H�E��E���E�����UH��AWSH��0��H�����I���     L�H�}�H��-     �    H��-     H�   H��-     H�H�E�H�E�   �    H��I��H��������H���H��-     H�  H��-     H�H�E�H�E�    �    H��I��H��������H���H�E�    �E�    ��   H�E������H�E�����H�E�H��H��H������   H!�H�E�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH�E��E��}��� �/���H��-     H�H�E��E�    ��   H�E�����H�E�����H�E�����H�E�H��H��H������   H!�H�E�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH�E�   H�E��E��}��  ����H��-     H�H�E�H��������H�H� H�� ����H��������H�H� H�� ����H��������H�H� H�� ����H�E�H��H��H��������H�H� H�� H������   H!�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH��������H�H� �����    H��0[A_]���UH��H�� ��H�����I���     L�H�}�u�H�E�H�E�H�E�� ����t�   �4�E�    �H�E�� ����t������H�E��E��E�9E�wڸ    ����UH��AWSH��0��H�����I��     Lۉ}̉u�H�U��}� u
�    �U  �H��-     ���u�H��-     ��PH��-     �H��-     H�H�E��E�    �E�    �E�    �  H�E�� ������  �U�H�E��H��H�T^������H��Ѕ��h  �E܉E��E�    �1  �    H��X������H���H�E�H�}� u'H�$�������H�<I�߸    H�u�������H�����H�E������}� tH�E������}� tH�E��P�����P��E�   H�E�H��H��H������   H!�H�E�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH�E��E��E�9E������I�߸    H�_P������H����H�E��E��}��� �L����}� t!�E���H�H�       H�H��H�E�H��H�E�H�     H��-     �    �E�H��0[A_]���UH��SH��H��H�����I���     L�H�}�H�}� �  H�E�H�E�H�E�H��%�  �E�H�E�H��%�  �E�H�E�H��%�  �E�H��������H�H� �U�Hc�H��H��P�����HH��H	��PH��H	��PH��H	��PH��H	��@��H��$H	�H��H������   H!�H��H�������  H!�H�EЋE�H�H��    H�E�H��P�����HH��H	��PH��H	��PH��H	��PH��H	��@��H��$H	�H��H������   H!�H��H�������  H!�H�EȋE�H�H��    H�E�H��@������  �H��-     ���u�H��-     ��PH��-     ��E�    �E�H�H��    H�E�H��P�����HH��H	��PH��H	��PH��H	��PH��H	��@��H��$H	�H��H������   H!�H�E�H�E�H��H��Y������H��ЋU�E��H�H��    H�E�H�������U�E��H�H��    H�E�H�������U�E��H�H��    H�E�H��P���P�P�� �P�P�� �P�P�� �P�P�� �P�P����P�U�E��H�H��    H�E�H��P���P�U�E��H�H��H��    H�E�H��@����t	�E������H��-     �    ����H��H[]���UH��H��8��H�����I�,�     L�H�}�H�U�H�����  �U�H�U�H�����  �U�H�U�H�����  �U�H��������H�H� �U�Hc�H��H��P�����HH��H	��PH��H	��PH��H	��PH��H	��@��H��$H	�H��H������   H!�H��H�������  H!�H�E�E�H�H��    H�E�H��P�����HH��H	��PH��H	��PH��H	��PH��H	��@��H��$H	�H��H������   H!�H��H�������  H!�H�E��E�H�H��    H�E�H��P�����HH��H	��PH��H	��PH��H	��PH��H	��@��H��$H	�H��H������   H!�H�E�H�E�����UH��SH����H�����I�Y�     L�H�}�H�E�H�E�H�E�L�@H�E�H�x�    ��Љ�H�U��2A��H�E�H���  �    H��[]���UH��SH����H�����I��     L�H�}�H�E�H�E�H�E�L�PH�E�L�HH�E�L�@�  ���މ�H�E��8A�2A�	A�H�E�L�PH�E�L�HH�E�L�@H�E�H�x�  ����A�A�1A��H�E�L�P H�E�L�H$H�E�L�@(H�E�H�x,�  ����A�A�1A���    H��[]���UH��SH����H�����I��     L؉}�H�u�H�U��E����H�E�0H�E���H��[]���UH��SH����H�����I�ɗ     L؉}�H�u�H�E�L�PH�E�L�HH�E�L�@�E���މ�H�E�8A�2A�	A�H�E� H��[]���UH��H����H�����I�a�     L؉}�H�u�H�U�E���2��H�E��H�E��    ����UH��H�� ��H�����I��     L؉}�u�U�H�E�    H�E�    �E��2H�E�H�U��E�H	E��E�H	E�H�E�H�U��M�0�    ����UH��AWSH����H�����I���     Lۉ}�I�߸    H��t������H��ҋE�� ����  ��H��    H��_ H�H��_ H�>��d   I��H��w������H����  H�0�������H�<I�߸    H�u�������H����  H�F�������H�<I�߸    H�u�������H����V  H�V�������H�<I�߸    H�u�������H����,  H�f�������H�<I�߸    H�u�������H����  �90  I��H��w������H�����   �90  I��H��w������H�����   �90  I��H��w������H����   �90  I��H��w������H����   �90  I��H��w������H����y�90  I��H��w������H����`�90  I��H��w������H����G�90  I��H��w������H����.�E�� ��H�v�������H�<I�߸    H�u�������H��Ґ�H��[A_]���UH��AWS��H�����I�g�     L�H� �������H��    �   �ƿ    I��H�70������H���H���������H��    �   �ƿ!   I��H�70������H���H�`�������H��    �   �ƿ"   I��H�70������H���H���������H��    �   �ƿ#   I��H�70������H���H�X�������H��    �   �ƿ$   I��H�70������H���H�P�������H��    �   �ƿ%   I��H�70������H���H���������H��    �   �ƿ&   I��H�70������H���H���������H��    �   �ƿ'   I��H�70������H���H���������H��    �   �ƿ(   I��H�70������H���H���������H��    �   �ƿ)   I��H�70������H���H�p�������H��    �   �ƿ*   I��H�70������H���H���������H��    �   �ƿ+   I��H�70������H���H���������H��    �   �ƿ,   I��H�70������H��А[A_]���UH��AWH����H�����I���     Lډ}�E��H���������H�<I�׸    H�u�������H��ѐH��A_]���UH��AWSH�� ��H�����I�a�     Lۉ}܃m�@I�߸    H��t������H��҃}�w8H�(      �E�H�H��H�E�U�H�E��H��I��H��������H����*�E܉�H��������H�<I�߸    H�u�������H��ҐH�� [A_]���UH��AWS��H�����I���     L�H�h�������H��    �   �ƿ@   I��H�70������H���H���������H��    �   �ƿA   I��H�70������H���H���������H��    �   �ƿB   I��H�70������H���H���������H��    �   �ƿC   I��H�70������H���H���������H��    �   �ƿD   I��H�70������H���H���������H��    �   �ƿE   I��H�70������H���H���������H��    �   �ƿF   I��H�70������H���H�8�������H��    �   �ƿG   I��H�70������H���H��������H��    �   �ƿH   I��H�70������H���H�X�������H��    �   �ƿI   I��H�70������H���H���������H��    �   �ƿJ   I��H�70������H���H���������H��    �   �ƿK   I��H�70������H���H���������H��    �   �ƿL   I��H�70������H���H���������H��    �   �ƿM   I��H�70������H���H���������H��    �   �ƿN   I��H�70������H���H���������H��    �   �ƿO   I��H�70������H���H�8�������H��    �   �ƿP   I��H�70������H���H��������H��    �   �ƿQ   I��H�70������H���H��������H��    �   �ƿR   I��H�70������H���H���������H��    �   �ƿS   I��H�70������H���H���������H��    �   �ƿT   I��H�70������H���H���������H��    �   �ƿU   I��H�70������H���H�(�������H��    �   �ƿV   I��H�70������H���H�H�������H��    �   �ƿW   I��H�70������H��А[A_]���UH��AWH����H�����I��     L�H�U�H�M�H�ο   I��H��h������H��ыE�H��A_]���UH��AWH��(��H�����I���     L؉}܋U܁� ������U��E�    �U�M�ο   I��H��h������H��Ѹ    H��(A_]���UH����H�����I�2�     L�H��     H�H�   �     �]���UH��AWSH����H�����I��     L�H�E�    �    H�ƿ  ��I��H��S������H���H�E�H��     H��   �    �   ��   �    �!   �(   ��   �   �!   �   ��   �   �!   �   ��   ��   �!   ��   ��   �H��     H�H�   � ����H��     H�H�   � %��� �E�M�H��     H�H�   H�E�H��     H�H�� �     H��     H�H���     H��     H�H   �    H��     H�H@  � !   H��     H�HP  � "' H��     H�H`  � # H��     H�Hp  � $  H��     H�H�   �   �    H�t������H��҉�H�[t������H��и    H�t������H��҉�H��������H�<I�߸    H�u�������H���H��     H�H��H��w������H��и    H��[A_]���UH��H����H�����I�l�     L؉}�H��     H�H�  H�E�������UH��H����H�����I�&�     L�H�}�H�E�H   �    H�E�H�  � 
   H�E�H�  � @� �    ����UH��H����H�����I�Ǉ     L�H��     H�H��   ��U�H��     H�H��   H�ыU��������H��     H�H���  �
   H��     H�H�  � 90  �����UH��H����H�����I�.�     L�H��     H�H��   ��U�H��     H�H   H�E�   ������UH��H����H�����I�̆     L�H�}��u�H�E��U�H�E�H��� ����UH��H����H�����I���     L�H�}��u�U�H�E��U�H�E�H��H�E�������UH��H����H�����I�B�     L؉}�H��-     H�H�U�H��-     �U�Hc�H�H�4�H��   H�4�H�U�H�U��U��Hc�H��    H�U�Hʋ�M���4	H��.     H�H��H�hy������H��и    ����UH��H����H�����I���     L؉}�H��-     H�H�U�H��-     �U�Hc�H�H�4�H������H�4�H�U�H�U��U��Hc�H��    H�U�Hʋ�M���4	H��.     H�H��H�hy������H��и    ����UH��SH��@��H�����I��     L�H�}��u܉�E��E��D�MD�E�} �u(�M0�U؈E�D�؈E�D�ЈE�D�ȈE�D���Eĉ��E����E��ȈE�H��-     H�H�E�H�E�H�E�H��-     �E�H�H��U؈��Eԃ���H��-     �E�H�H��Ƀ�H��H��H���H	�H���EЃ���H��-     �E�H�H��Ƀ�H��H��H���H	�H���Ẽ���H��-     �E�H�H��Ƀ�H��H��H���H	�H���Eȃ���H��-     �E�H�H��Ƀ�H��H��H���H	�H���Eă���H��-     �E�H�H��Ƀ�H��H��H��H	�H���E�����H��-     �E�H�H��Ƀ�H��H��H��H	�H���E�����H��-     �E�H�H��Ƀ�H��H��H��H������H	�H��H��-     �E�H�H��H�H�H�P�E���E��H�H��    H�E�HЋ�E܃�� H�E���H��H�hy������H��ЋE��H�H��H��    H�E�HЋ�E܃���HH�E���H��H�hy������H��и    H��@[]���UH��SH����H�����I��     L�H�}��E�    �F�E��@�Ћu�H�E�j jj j j A�    A�    �    H��H�{������H���H��(�E��}�~��    H�]�����UH��AWSH����H�����I���     L�H�E�    �   H�ƿ  ��I��H��S������H���H�E�H��.     H�H��.     H��    �    H��H�hy������H���H��.     H�H��H��}������H��и    H��[A_]���UH��AWH����H�����I�Հ     L؉}�}� t3�U�Hc�Hi�gfffH�� ����)щ�Hc�H��I��H���������H��ҐH��A_]���UH��AWATSH����H�����I�g�     L�H�@/     H�    H��.     H���������H�H�H� /     H��   �    I��H��^������H���H� /     H�H��.     H�H��.     H��p  �    H��I��H��������H���H�@/     H�H�PH�@/     H�H��.     H�H���   H��.     H�H`  H��I��H�4������H���H��.     H�Hǀ�      H��.     H�Hǀ�      H��.     H�Hǀ�     H��������H�H�H��.     H�H���   H��.     L�$H�-�������H�4�    I��H���������H���I��$�   H��.     L�$H�3�������H�4�    I��H���������H���I��$�   H��.     L�$H�:�������H�4�    I��H���������H���I��$   H��.     L�$H�A�������H�4�    I��H���������H���I��$  H��.     L�$�   I��H�R�������H���I��$  H��.     H�Hǀ�       H��.     H�Hǀ`      H��.     H�H��.     H�H��.     H�H��.     H�H��.     H�H���   H��[A\A_]���UH��AWATSH��h��H�����I�+}     L�H�}�H�u�H�U�H�M�D�E�D�M�H�E�H�¾   �    I��H��^������H���H�E��p  �    H��I��H��������H���H�@/     H�H�PH�@/     H�H�U�H���   H�E�H`  H��I��H�4������H���H�E�H�U�H�P8H�E�H�U�H�P@�E�������   H�E�Hǀ�      H�E�Hǀ�   #   H�E�H�¾   �   I��H��^������H���H�E��  �    H��I��H��������H���H�E�H�U�H��P  H�E�Hǀ�      H�E�Hǀ�   2  �F�E�����u<H�E�Hǀ�      H�E�Hǀ�      H�E�Hǀ�       H�E�Hǀ�     �E�%�   ��tH�E�H���   H�E��ʀH���   H�E�H�U�H���   L�e�H�-�������H�4�    I��H���������H���I��$�   L�e�H�3�������H�4�    I��H���������H���I��$�   L�e�H�:�������H�4�    I��H���������H���I��$   L�e�H�A�������H�4�    I��H���������H���I��$  L�e��   I��H�R�������H���I��$  H�E�H���   H�E�H�� H���   �E�������   H�E�H�¾   �   I��H��^������H���H�E�H�U�H��  H�E�H���   H�E�H��H���   H�E�H�E�H�Eк   �    H��I��H��������H���H��������H��PH�EЉPH��������H��PH�EЉPH��������H��PH�EЉPH��������H��PH�EЉPH�E�H���������H�H�H��   H�E�H���   H�E�H�PH�E�H���   H�E�H�PH�E�H��   H�E�H�P(H�U�H�E�H��  H�P H�E�H�U�H�PH�E�H�@H    H�U�H�E�H��P  H�PPH�E�H��  H�E�H�PXH�E�H��  H�E�H�H�E��U�Hc�H�P`H�E�H�UH�PhH�E�H�UH�PpH�E�Hǀ`      H� /     H�H�E��H�E�H��`  H�E�H�E�H��`  H��u�H�U�H�E�H��`  H�E�H��h[A\A_]���UH��AWSH��P��H�����I�x     L�H�}�H�u�H�U�H�M�D�E�D�M�H�E H�E�H�E�H�¾   �    I��H��^������H���H�Eغp  �    H��I��H��������H���H�@/     H�H�PH�@/     H�H�U�H���   H�E�H`  H��I��H�4������H���H�E�H�U�H�P8H�E�H�U�H�P@�E�������   H�E�Hǀ�      H�E�Hǀ�   #   H�E�H�¾   �   I��H��^������H���H�Eк  �    H��I��H��������H���H�E�H�U�H��P  H�E�Hǀ�      H�E�Hǀ�   2  �F�E�����u<H�E�Hǀ�      H�E�Hǀ�      H�E�Hǀ�       H�E�Hǀ�     H�E�H�U�H���   H�E�H�U�H���   H���   H�E�H�U�H���   H���   H�E�H�U�H��   H��   H�E�H�U�H��  H��  H�E�H�U�H��  H��  H�E�H�U�H��  H��  H�E�H���   H�E�H�PH�E�H���   H�E�H�PH�E�H��   H�E�H�P(H�U�H�E�H��  H�P H�E�H�U�H�PH�E�H�@H    H�U�H�E�H��P  H�PPH�E�H��  H�E�H�PXH�E�H��  H�E�H�H�E؋U�Hc�H�P`H�E�H�UH�PhH�E�H�UH�PpH�E�Hǀ`      H� /     H�H�E��H�E�H��`  H�E�H�E�H��`  H��u�H�U�H�E�H��`  H�U�H�E�H��h  H�E�H��P[A_]���UH��H����H�����I�pt     L�H� /     H�H�U��#H��.     H�H9U�tH�U�H��`  H�U�H�}� u���H�}� �  H��.     H�H��.     H�H��.     H�H��.     H�H�
H��.     H�H�x/     H�H�JH��.     H�H��.     H�H�JH��.     H�H��.     H�H�JH��.     H�H��/     H�H�J H��.     H�H��.     H�H�J(H��.     H�H� /     H�H�J0H��.     H�H�/     H�H�J8H��.     H�H�h/     H�H�J@H��.     H�H�(/     H�H�JHH��.     H�H��.     H�H�JPH��.     H�H�`/     H�H�JXH��.     H�H�P/     H�H�J`H��.     H�H��.     H�H�JhH��.     H�H�X/     H�H�JpH��.     H�H��/     H�H�JxH��.     H�H�0/     H�H���   H��.     H�H��.     H�H���   H��.     H�H��.     H�H���   H��.     H�H��/     H�H���   H��.     H�H�/     H�H���   H��.     H�H�H/     H�H���   H��.     H�H�8/     H�H���   H��.     H�H��.     H�H���   H��.     H�H�/     H�H���   �E�    �:H��.     H��U�Hc�H�H��.     H��2�U�Hc�@��`  �E��}��  ~�H��.     H�H��`  H��.     H�H��.     H�H���   ��   H��uH��.     H�H���   H��u#H��.     H�H��`  H��.     H�H��.     H�H��uH� /     H�H��.     H�H��.     H�H��.     H�H��.     H�H�H��.     H�H��.     H�H�RH�x/     H�H��.     H�H�RH��.     H�H��.     H�H�RH��.     H�H��.     H�H�R H��/     H�H��.     H�H�R(H��.     H�H��.     H�H�R0H� /     H�H��.     H�H�R8H�/     H�H��.     H�H�R@H�h/     H�H��.     H�H�RHH�(/     H�H��.     H�H�RPH��.     H�H��.     H�H�RXH�`/     H�H��.     H�H�R`H�P/     H�H��.     H�H�RhH��.     H�H��.     H�H�RpH�X/     H�H��.     H�H�RxH��/     H�H��.     H�H���   H�0/     H�H��.     H�H���   H��.     H�H��.     H�H���   H��.     H�H��.     H�H���   H��/     H�H��.     H�H���   H�/     H�H��.     H�H���   H�H/     H�H��.     H�H���   H�8/     H�H��.     H�H���   H��.     H�H��.     H�H���   H�/     H�H��.     H�H���   H�p/     H��E�    �9H��.     H�H��.     H�4�U�Hc�H֋U�Hc���`  ��E��}��  ~�������UH��H����H�����I��k     L�H� /     H�H�U��#H��.     H�H9U�tH�U�H��`  H�U�H�}� u���H�}� �
  H�U�H���   ��   H���B  H��.     H�H�U�H�
H�x/     H�H�U�H�JH��.     H�H�U�H�JH��.     H�H�U�H�JH��/     H�H�U�H�J H��.     H�H�U�H�J(H� /     H�H�U�H�J0H�/     H�H�U�H�J8H�h/     H�H�U�H�J@H�(/     H�H�U�H�JHH��.     H�H�U�H�JPH�`/     H�H�U�H�JXH�P/     H�H�U�H�J`H��.     H�H�U�H�JhH�X/     H�H�U�H�JpH��/     H�H�U�H�JxH�0/     H�H�U�H���   H��.     H�H�U�H���   H��.     H�H�U�H���   H��/     H�H�U�H���   H�/     H�H�U�H���   H�H/     H�H�U�H���   H�8/     H�H�U�H���   H��.     H�H�U�H���   H�/     H�H�U�H���   �S����%H�U�H���   ��   H��uH�U�H��`  H�U�H�}� u���H�}� �p  H��.     H�U�H�H�U�H�H��.     H�H�U�H�RH�x/     H�H�U�H�RH��.     H�H�U�H�RH��.     H�H�U�H�R H��/     H�H�U�H�R(H��.     H�H�U�H�R0H� /     H�H�U�H�R8H�/     H�H�U�H�R@H�h/     H�H�U�H�RHH�(/     H�H�U�H�RPH��.     H�H�U�H�RXH�`/     H�H�U�H�R`H�P/     H�H�U�H�RhH��.     H�H�U�H�RpH�X/     H�H�U�H�RxH��/     H�H�U�H���   H�0/     H�H�U�H���   H��.     H�H�U�H���   H��.     H�H�U�H���   H��/     H�H�U�H���   H�/     H�H�U�H���   H�H/     H�H�U�H���   H�8/     H�H�U�H���   H��.     H�H�U�H���   H�/     H�H�U�H���   H�p/     H���������UH��H����H�����I�ef     L�H�}�H� /     H�H�E��&H�E�H���   H9E�uH�E��H�E�H��`  H�E�H�}� uӸ    ����UH��AWSH���   ��H�����I��e     Lۉ�,���H�� ���H�����H������E�    �@   I��H�R�������H���H�E�H������    �   H��I��H���������H����E�    �   H�����H�E�H�Ѻ   �   H��I��H���������H���H�E��   H��H�F�������H�<I��H�G�������H��Ѕ�u4H�E�H�xH�����H���8   �   I��H���������H��ЃE���E��}��  �^����}� u#H�E�H��I��H���������H��и    �	  H�E�H�@(��H�E�H�@)�  �E��E����  ��H����E�E�%�  ��t�E��E䍐�  ��H���	�E��E�%�  ��t�E�HǅP���    HǅH���    Hǅ@���    Hǅ8���    H��P���H�¾   �    I��H��^������H���H��P����   �    H��I��H��������H���H��H���H�¾   �    I��H��^������H���H��H����   �    H��I��H��������H���H��@���H�¾   �    I��H��^������H���H��@����   �    H��I��H��������H��ЋE�H��8����ƿ    I��H��^������H��ЋE�H�����H��8����    H��I��H��������H���H��������H�H�H��P����   H��H��I��H�o�������H���H��8���H�E��E�    ��   I�߸    H��X������H���H��X���H�E�����H�E�����H�E�����H��X���H��H��H������   H!�H�E�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH�E��E��E�;E�����H��@���H�E�H��8���H�E��E�    ��   H�E�H��I��H��d������H���H�E�H�E�����H�E�����H�E�����H�E�H��H��H������   H!�H�E�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH�E�   H�E��E��E�;E������H��@���H��I��H��d������H���H�E�H��H�������H��H�������H��H�������H�E�H��H��H��H���H������   H!�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH��H���H��I��H��d������H���H�E�H��P���H������H��P���H������H��P���H������H�E�H��H��H��P���H��H������   H!�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH��P���H��I��H��d������H���H�E� �H�E�H�E�H��I��H��P������H����E��   ��m��}� �H������   �    H��I��H���������H���H�����H��I��H�c�������H��ЉE�H�����H��I��H��������H��ЋE����¾    H�    �   I��H��������H��ЋE�H�����H�щ¾   H�    �   I��H���������H��ЋE�H�H�  ��   H�H��x���H��x���H��p���H��x���   H��x���H��h���H��x���   �E�    �1�E���Hc�H��x���HE�H�H��    H��h���H�H��E��}�~�H����� t&H�����H��p���H��H��I��H��������H���H�� ��� td�E�    �P�E�H�H��    H�� ���H�H��E�H�H��    H��h���H�H� H��H��I��H��������H��ЃE��E�;�,���|�H�E�H��I��H��P������H����E��   ��m��}� �H���������H�H� H���E�H�H�    �   H�H��H�E�H�@H�ǋ�,���H�E���p�����h���A��A�   H��I��H�Ă������H���H��H��`���H��P���H��H��`���H��(  H��H���H��H��`���H��0  H��@���H��H��`���H��8  H��8���H��H��`���H��@  �E�Hc�H��`���H��H  H�E�H��I��H���������H���H��`���H���   H�e�[A_]���UH��AWSH���   ��H�����I��Z     Lۉ�,���H�� ���H�����H�����L������E�    �@   I��H�R�������H���H�E�H������    �   H��I��H���������H����E�    �   H�����H�E�H�Ѻ   �   H��I��H���������H���H�E��   H��H�F�������H�<I��H�G�������H��Ѕ�u4H�E�H�xH�����H���8   �   I��H���������H��ЃE���E��}��  �^����}� u#H�E�H��I��H���������H��и    �	  H�E�H�@(��H�E�H�@)�  �E��E����  ��H����E�E�%�  ��t�E��E䍐�  ��H���	�E��E�%�  ��t�E�HǅP���    HǅH���    Hǅ@���    Hǅ8���    H��P���H�¾   �    I��H��^������H���H��P����   �    H��I��H��������H���H��H���H�¾   �    I��H��^������H���H��H����   �    H��I��H��������H���H��@���H�¾   �    I��H��^������H���H��@����   �    H��I��H��������H��ЋE�H��8����ƿ    I��H��^������H��ЋE�H�����H��8����    H��I��H��������H���H��������H�H�H��P����   H��H��I��H�o�������H���H��8���H�E��E�    ��   I�߸    H��X������H���H��X���H�E�����H�E�����H�E�����H��X���H��H��H������   H!�H�E�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH�E��E��E�;E�����H��@���H�E�H��8���H�E��E�    ��   H�E�H��I��H��d������H���H�E�H�E�����H�E�����H�E�����H�E�H��H��H������   H!�H�E�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH�E�   H�E��E��E�;E������H��@���H��I��H��d������H���H�E�H��H�������H��H�������H��H�������H�E�H��H��H��H���H������   H!�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH��H���H��I��H��d������H���H�E�H��P���H������H��P���H������H��P���H������H�E�H��H��H��P���H��H������   H!�H�у������H��	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��H�����H�� 	�HH��$���у��P���	ʈPH��P���H��I��H��d������H���H�E� �H�E�H�E�H��I��H��P������H����E��   ��m��}� �H������   �    H��I��H���������H���H�����H��I��H�c�������H��ЉE�H�����H��I��H��������H��ЋE����¾    H�    �   I��H��������H��ЋE�H�����H�щ¾   H�    �   I��H���������H��ЋE�H�H�  ��   H�H��x���H��x���H��p���H��x���   H��x���H��h���H��x���   �E�    �1�E���Hc�H��x���HE�H�H��    H��h���H�H��E��}�~�H����� t&H�����H��p���H��H��I��H��������H���H�� ��� td�E�    �P�E�H�H��    H�� ���H�H��E�H�H��    H��h���H�H� H��H��I��H��������H��ЃE��E�;�,���|�H�E�H��I��H��P������H����E��   ��m��}� �H���������H�H� H���E�H�H�    �   H�H��H�E�H�@H�ǋ�,���H�E�H���������p�����h���A��A�   H��I��H��������H���H�� H��`���H��P���H��H��`���H��(  H��H���H��H��`���H��0  H��@���H��H��`���H��8  H��8���H��H��`���H��@  �E�Hc�H��`���H��H  H�E�H��I��H���������H���H��`���H���   H�e�[A_]���UH��AWH��(��L�����I��O     M�H�}�H�u�H�U�H�M�H�E�H��H�O�������I�< M�Ǹ    H�u�������L��ҐH��(A_]���UH��AWH��(��H�����I�iO     L�H�}�H�u�H�U�H�M�H�U�H��I��H��������H��ҐH��(A_]���UH��AWH��(��H�����I�O     L�H�}�H�u�H�U�H�M�H�U�H��I��H�<m������H��ҐH��(A_]���UH��H�� ��H�����I��N     L�H�}�H�u�H�U�H�M�H�M�H���������H�H�
H���������H�H�H��  H�X�������H�H������UH��AWSH��0��H�����I�CN     L�H�}�H�u�H�U�H�M�H�E�    H�E���H�E�H�ο   I��H��^������H���H�E�H��/     H��H��0[A_]���UH��AWH��(��H�����I��M     L�H�}�H�u�H�U�H�M�H�U�H��I��H�qa������H��ҐH��(A_]���UH��AWSH�� ��H�����I�jM     L�H�}�H�u�H�U�H�M�H�U�H�EЉ�H�E�H��H�¿    I��H�5<������H���H�H��/     H��H�� [A_]���UH��AWSH�� ��H�����I��L     L�H�}�H�u�H�U�H�M�H�U�H�EЉ�H�E�H��H�¿    I��H�K=������H���H�H��/     H��H�� [A_]���UH��AWSH��0��H�����I�rL     L�H�}�H�u�H�U�H�M�L�E�H��������H�H�U�H�H��������H�H�U�H�PH��������H�H�U�H�PH��������H�H�U�H�PH���������H�H� H���   H��������H�H�P H�}� tcH�}�tH�}�uUH�U�H���������H�H� H��H��I��H��������H���H���������H�H� H��H��������H�H�P(�H��������H�H�@(    ��H��0[A_]���UH��AWSH��@��H�����I�+K     L�H�}�H�E�H�E�H�E�H�PH�U�� tH�E�H�PH�U�� mH�E�H�PH�U�� pH�E��  H���������H�� �HH���������H��
H�U�H�։�I��H�w�������H���H��H�E�H��H��I��H��������H��АH��@[A_]���UH��AWH��H��H�����I�^J     L�H�}�H�u�H�U�H�M�L�E�L�M�H�UȉU�H�}�	v�E�    H��      �U�Hc�H�H��H�U�L�M�L�E�H�M�H�U�H�u�H�}�H���u�I��I��������I�A��H���L�}�����UH��AWH����H�����I��I     L�H��������H���A�    �   �   �r   I��I��0������I�A�ѐH��A_]�f���AWAVAUATASARAQAPWVUTSRQP�%�A H�L$H�T$H�t$0H�|$8L�D$@�����%�A XYZ[\]^_AXAYAZA[A\A]A^A_��H�%0#E H��   H�h    hr   �z�����UH��AWSH��  ��H�����I��H     L��E�    �E� H�������   �    H��I��H��������H���H���������H�<I�߸    H�u�������H���H�(�������H�H� H��I��H�"�������H��ЈE�}� ��  ��E��H��������H�<I�߸    H�u�������H��Ҹ    �怀}�
�d  �}� ��   �E�    ��   H�H      �E�Hc�H�H��H�H�H��H�H�H������H��H��I��H���������H��Ѕ�u\H�H      �E�Hc�H��H�H�H��H�H�H��H� H��H��     H�H��     H�H������H�ƿ   ���L�}�u8�H������H��H��������H�<I�߸    H�u�������H��Ҹ    �怃E��}�����H�������   �    H��I��H��������H����E�    �H��������H�<I�߸    H�u�������H��Ҹ    ���M�}�u�}� ~�m��E�H�Ƅ���� �.�}�u�E�H��U爔������E�P�U�H��U爔������������UH��AWH����H�����I�F     L؉}�H�u��H�!�������H�<I��H��������H��Ҹ    �怸    H��A_]���UH��AWH����H�����I��E     L؉}�H�u��H�!�������H�<I��H��������H��Ҹ    �怸    H��A_]���UH��AWH����H�����I�VE     Lډ}�H�u��I�׸    H���������H��Ѹ    �怸    H��A_]���UH��AWH����H�����I��D     L؉}�H�u��H�!�������H�<I��H��������H��Ҹ    �怸    H��A_]���UH��AWH����H�����I��D     Lډ}�H�u��I�׸    H�K�������H��Ѹ    �怸    H��A_]���UH��AWH����H�����I�?D     L؉}�H�u��H�!�������H�<I��H��������H��Ҹ    �怸    H��A_]���UH��AWH����H�����I��C     L؉}�H�u��H�!�������H�<I��H��������H��Ҹ    �怸    H��A_]���UH��AWSH��   ��H�����I�uC     Lۉ�l���H��`���H��p�����   �    H��I��H��������H���H��p���H��I��H�g������H����H��p���H��H�@�������H�<I�߸    H�u�������H��Ҿ   �    I��H���������H��и    �怸    H�Đ   [A_]���UH��AWSH�� ��H�����I��B     Lۉ}�H�u��H�r�������H�<I��H��������H����E�    ��   H�H      �E�Hc�H�H��H�H�H��H�H� H��I��H��������H���H�H      �E�Hc�H�H��H�H�H��H�H� H��I��H�a�������H��ЉE���    I��H���������H��ЃE��}�~�H�H      �E�Hc�H�H��H�H�H��H�H��H� H��I��H��������H��п
   I��H���������H��ЃE��}�� ����    �怸    H�� [A_]���UH��AWH����H�����I�*A     L؉}�H�u��H�!�������H�<I��H��������H��Ҹ    �怸    H��A_]���UH��AWH����H�����I��@     L؉}�H�u��H�!�������H�<I��H��������H��Ҹ    �怸    H��A_]���UH��AWH����H�����I�d@     L؉}�H�u��H�!�������H�<I��H��������H��Ҹ    �怸    H��A_]���UH��AWH����H�����I�@     L؉}�H�u��H�!�������H�<I��H��������H��Ҹ    �怸    H��A_]���UH��AWH����H�����I��?     L؉}�H�u��H�!�������H�<I��H��������H��Ҹ    �怸    H��A_]���UH��AWH����H�����I�;?     L؉}�H�u��H�!�������H�<I��H��������H��Ҹ    �怸    H��A_]���UH��AWH����H�����I��>     Lډ}�H�u��I�׸    H��h������H��Ѹ    �怸    H��A_]���UH��AWH����H�����I�~>     L؉}�H�u��H�!�������H�<I��H��������H��Ҹ    �怸    H��A_]���UH��AWSH�� ��H�����I�>     L�H�}�H�E�H��P  H�E��E�    �=H�E�@��u(H�E�H� H��tH�E�H� H��I��H�qa������H���H�E��E��}��   ~�H�E�H��I��H�qa������H��АH�� [A_]���UH��AWSH��P��H�����I�n=     Lۉ}�H�u�H�E�H�E��H�E�Hǀ�      H�E�H��h  H�E�H�}� u�H�E�    H�E�    f�E�H�E�H��  H�E�H��H��I��H�)�������H���H�E�H�E��  H�E�H��@  H�E��E�    �H�E��P�����HH��H	��PH��H	��PH��H	��PH��H	��@��H��$H	�H��H������   H!�H�E�H�E�H��I��H��Y������H���H�E��E��E�Hc�H�E�H��H  H9��g���H�E�H��(  H��I��H�qa������H���H�E�H��0  H��I��H�qa������H���H�E�H��8  H��I��H�qa������H���H�E�H��@  H��I��H�qa������H���H�E�H��H���������H���H�E�H���   �� H����   H�E�H���   H��I��H�Ô������H���H�E�H���   H��I��H�Ô������H���H�E�H��   H��I��H�Ô������H���H�E�H��  H��I��H�Ô������H���H�E�H��  H��I��H���������H���H�E�H��h  H�E�H�}� �����H�p�������H��  H�E�H�E��   H�E�H�E�H�@�������H�H� H�E��8H�E�H��`  H9E�uH�E�H��`  H�E�H��`  �H�E�H��`  H�E�H�}� u�H�E�H��h  H�E�H�E�H��I��H�qa������H���H�}� �o���H�p�������H�� �H��P[A_]���UH��H����H�����I��9     L؉�f�E��m������UH��H����H�����I��9     L��E�#  �U��E�����UH��H����H�����I��9     L؉}��]������UH��H����H�����I�U9     L�H�}��E������UH��H����H�����I�&9     L�H�}��M������UH��AWSH����H�����I��8     L�H�U�H�E�H�ƿ   I��H��g������H��ЋE�%   ��u"H�}�������H�<I��H��������H�����H���������H�<I��H��������H��� �   "� �f���f��"���I�߸    H�)������H��Ҹ    H��[A_]���UH��H�� ��H�����I� 8     L؉}�u�U�M��E���%  � �E���% � 	E���%   	E�%�   	�   ���  ��  ���E��E�����UH��H����H�����I��7     L؉}��u��U�M�D�E�E���%  � �E���% � 	E���%   	E�%�   	�   ���  �E��  �����UH��H�� ��H�����I�(7     L؉}�u�U�M��E���%  � �E���% � 	E���%   	E�%�   	�   ���  ��  ���E��E�����UH��H����H�����I��6     L؉}��u��U�M�D�E�E���%  � �E���% � 	E���%   	E�%�   	�   ���  �E��  �����UH��AWSH��0��H�����I�-6     L�H�}ȉu��E�����H� �������H�<I�߸    H�u�������H����E�    �  �E�    �h  �E�    �N  �U�u�E�   ��H���������H��ЉE܃}���  �E�    ��   H�      �E�Hc�H�H��H�H�H��Hȋ %��� �E���9�t	�E��   H�      �E�Hc�H�H��H�H�H��H�H�@H��H��������H�<I�߸    H�u�������H��ҋM�U�E��H��������H�<I�߸    I�u�������I�A����}��   �2����}�   u:�u�M�U�E�A����H�(�������H�<I�߸    I�u�������I�A�����E��}�������E��}�������E��E�;E��r����    H��0[A_]���UH��H��(��H�����I�.4     L؉}��E������E�    �   �E�    �~�E�    �k�E���%  � �E���% � 	E���%   	�  ���  ��  ���E�E�E��E���9E�u�E���    �E�E�����.�E��}�~��E��}��x����E��}��   �^������������UH��H��(��H�����I�K3     L؉}��E������E�    �E�    �   �E�    �   �E�    �o�E���%  � �E���% � 	E���%   	�  ���  ��  ���E�E�E��E����E�9�u�E���E�U���	ЉE�E��.�E��}�v��E��}��t����E��}��   �W������������UH��H��(��H�����I�Z2     L؉}܉u��E������E�    �E�    �   �E�    �   �E�    �y�E���%  � �E���% � 	E���%   	�  ���  ��  ���E�E�E��E���9E�u'�E�����9E�u�E���E�U���	ЉE�E��.�E��}�~��E��}��j����E��}��   �M������������UH��H��0��H�����I�\1     L؉}܉u؉U��E������E�    �   �E�    �   �E�    �   �E���%  � �E���% � 	E���%   	�  ���  ��  ���E�E�E��E���9E�u5�E�����9E�u'�E�����9E�u�E���E�U���	ЉE�E��2�E��}��o����E��}��U����E��}��   �8������������UH��H����H�����I�M0     L؉�f�E��    ����UH��H����H�����I�0     L؉}��u��U��f�E�    ����UH��H����H�����I��/     L؉}�u�E�#E�E��E���!E��E�����UH��AWSH��@��H�����I��/     Lۉ}��u��U��U��u��E��    ��I��H���������H��ЉE�E�����H��/     f��E��H��/     f�T�U��u��E��   ��I��H���������H��Љ�H�E��U��u��E��   ��I��H���������H��Љ�H�E؋U��u��E��   ��I��H���������H��Љ�H�EЋU��u��E��   ��I��H���������H��Љ�H�EȋU��u��E��    ��I��H���������H��Љ�H�E�H�E�H�� HE�H���H��H��/     H�TH�E�H�� HE�H���H��H��/     H�TH�E����H��/     H�D�    H��@[A_]���UH��AWSH����H�����I��-     Lۺ8   �    H��/     H�<I��H��������H��п   I��H���������H��ЉE�}��u/H�X�������H�<I�߸    H�u�������H��Ҹ������   H���������H�<I�߸    H�u�������H��ҋE��ЋE������M����Ɖ�H�R�������H���H��/     �D��H��/     �����H���������H�<I�߸    H�u�������H���H��������H��@ ��H�E�    �  � H��I��H��S������H���H�U�H��������H�H�P0�   H��[A_]���UH��H��8��H�����I�a,     L�H�}�H�u�H�U�H�E�6  H�E�H��� ����H�U�H�����������   	ЉE�H�E�H��� ����H�U�H�����������   	ЉE��E�    �,  H�E�H�P�E���H�H�H   H�E��E�H�H��H��H�E�HE��E�H�H��H��H�E�HE�B�E�H�H��H��H�E�HЋ�E�H�H��H��H�E�H����P�E����E�H�H��H��H�E�HȉP�U�H�Eȉ�U�H�EȉPH�E��@    �E�H�H��H��H�E�HЋ@��?��t5�E�H�H��H��H�E�HЋ@����H�EȉH�Eȋ ������H�Eȉ�E�H�H��H��H�E�HЋ ��f%���H�E�������� 	�f���҃��у��P���	ʈP�E�H�H��H��H�E�HЋ@��f%���H�E������H�� 	�Hf���҃��у��P���	ʈPH�Eȋ ��f%���H�E������H�� 	�Hf���҃��у��P���	ʈPH�Eȋ@��f%���H�E������H�� 	�Hf���҃��у��P���	ʈP�E��}������������UH��H����H�����I��)     L�H�}�H�E�H�@H  �H�E�H�@H  H����%����H�E�H�@H  �H�E�H�@H  H���Ѐ�������UH��H����H�����I�)     L�H�}�H�E�H�@H  �H�E�H�@H  H����   ��H�E�H�@H  �H�E�H�@H  H���Ѐ�������UH��H����H�����I��(     L�H�}�H�E�H�@H� �H�E�H�@H� H����%����H�E�H�@H� �H�E�H�@H� H����%���������UH��H����H�����I�
(     L�H�}�H�E�H�@H� �H�E�H�@H� H����   ��H�E�H�@H� �H�E�H�@H� H����   �������UH��H����H�����I��'     L�H�}�H�E�H�@H  �H�E�H�@H  H����%���?�H�E�H�@H �H�E�H�@H H����%���?������UH��H����H�����I�'     L�H�}�H�E�H�@H  �H�E�H�@H  H����   ��H�E�H�@H �H�E�H�@H H����   �������UH��H����H�����I��&     L�H�}������UH��H����H�����I�b&     L�H�}�H�E�H�@H`  �  ������UH��H����H�����I�#&     L�H�}��  ���E��E��� �E��E���  �H�E�H�@H  �H�E�H�@H  H����   ��H�E�H�@H  �H�E�H�@H  H����%�����H�E�H�@H  �H�E�H�@H  H����   �������UH��H����H�����I�[%     L�H�}������UH��H����H�����I�0%     L�H�}�H�E�H�@HQ  �    H�����UH��H����H�����I��$     L�H�}��H�E�H�@HQ  � %   ��t琐����UH��SH��8��H�����I��$     L�H�}Љu�H�U��M��E�    �E�    H�E�H�E��E���%  ��E����	�  F�E�H�E�H��H���������H���H�E�H�@H Q  H�E��H�E�H�@HQ  H�E��E�    �   H�E�H��H��������H���H�E�H�@HQ  � �E܋E�Hc�H�E�HЋU܈�E��9E�~�E������E�H�H�PH�E�HЉʈ�E��9E�~�E������E�H�H�PH�E�HЉʈ�E��9E�~�E������E�H�H�PH�E�HЉʈ�E��E�;E��?���H�E�H��H���������H��АH��8[]���UH��H����H�����I�#     L؉}�H�u��U������UH��H��8��H�����I��"     L؉}�H�u�H�U�H�E�H�E��E�    �   �E���H�H��    H�E�H�H�E��E�    �k�U��������E��Hc�H�E�H�� ���E�}�u�E�H�H��    H�E�HE܉� �}�u�E�H�H��    H�E�H��  ��E��}�~��E��}��]���������UH��SH����H�����I��!     L�H�}��E�    �H�E�H�P,�E���H�H��     �E��}��  ~�H�E�H�@,H��H���������H�H�ο����H��������H���H��������H��@��E�H��������H��@��E�H�E�H�@H�  �    �E�%�  �E���%  �	�H�E�H�@H�  �H�E�H�@H�  �   p �H��[]���UH��H����H�����I��      L؉}��u�H���������H��R4��t7�U��с��  �U�����  �	�H���������H�H�@H�  �ʉ������UH��H����H�����I�t      L�H�}�H�(0     H�H�M�H)�H�`0     H�H�����UH��AWSH��@��H�����I�!      L�H�}�H�E�H�h0     H��E� H�E�H�E��E�    �H�E�� ���E�ЈE�H�E��E��}�~߀}� t/H���������H�<I�߸    H�u�������H��Ҹ   �4  H�h0     H�H��H�EӺ   H��H��I��H�o�������H���H�h0     H�H�H	H�E̺   H��H��I��H�o�������H����E� �E� H�h0     H��@��%  ��H�(0     H�H�(0     H��    �  @ H�`0     H�43H��I��H��S������H���H�h0     H��@<��   H���������H�<I�߸    H�u�������H���H�h0     H��@��H��H���������H���H��H�H0     H�H�h0     H�H�@H��H���������H���H��H�@0     H��   H�h0     H��@��unH���������H�<I�߸    H�u�������H���H�h0     H��@��H��H���������H���H��H�H0     H�H�@0     H�    H�E�H��H��������H�<I�߸    H�u�������H��Ҹ    H��@[A_]���UH��H�� ��H�����I�?     L�H�}�H�u�H�E� �E�H�E�� �E��E�;E�u�    ����������UH��SH��8��H�����I��     L�H�}�H�u�H�U�H�H0     H�H��$H�E�H�E�H�E�H�H0     H��@��$�E��E�    �SH�E�H�PH�U�� ��H��H���������H���H�E�H�E�H�U�H��H��H���������H��Ѕ�uH�E���E��E�;E�|��    H��8[]���UH��AWSH����H�����I�     L�H� 0     H��@@��f�f�E��E��������*  H� 0     H��@0���
  H� 0     H��@4����   H� 0     H��@4H� 0     H��R0��E�    �CH� 0     H��@@��f�f�E��E�������t#����I��H��&������H��ЃE��}�	~���H� 0     H��@D��tN�CH� 0     H��@D��f�f�E��E�������t#����I��H��&������H��ЃE��}�	~����}�	�    ��������������    H��[A_]���UH��H��0��H�����I��     L�H�E�   H�E�H   H�E�  � ���E��e��&H�E�H� H�E�H�RSD PTR H9E�uH�E��[H�E�H�E�H;E�rЋE�H�E�H�E�H   H�E��&H�E�H� H�E�H�RSD PTR H9E�uH�E��H�E�H�E�H;E�rи    ����UH��AWSH�� ��H�����I��     L�H��������H�<I�߸    H�u�������H��Ҹ    H�i�������H���H�E�H�}� ��   H�E�H��H���������H���H�@0     H�H�H0     H�H�0�������H�H��H��H�	�������H���H��H� 0     H�H� 0     H��@(��H��H���������H���H�E�H�E�H�P0     H�H�E�H�A�������H�4H��H���������H��Ѕ��!  �*H�5�������H�<I�߸    H�u�������H����  H�P0     H�H��$H�E�H�P0     H��@�E��   H�E�   H�F�������H�4H��I��H�G�������H��Ѕ�u~H�E�H�E�� ����H���H��HE�H�E�� <
uH�E�H�E�� f���
��H�00     f�H�E�H�E�� <
uH�E�H�E�� f���
��H�X0     f��=H�E��E�P��U���<����%H�K�������H�<I�߸    H�u�������H���H�� [A_]���UH����H�����I�3     L�H�00     ��� ��H� 0     H��R@f�H� 0     H��@D��t'H�X0     ��� ��H� 0     H��RDf�]���UH��AWH����H�����I��     L��H�h0     H��@<v(H� 0     H����   H� 0     H�H�Rx�H�`�������H�<I�ϸ    H�u�������H����E���d   ���E��E�E��E����u��   �d   ������UH��H�� ��H�����I��     L�H�}�u�H� �Ƥ~� H�E��E�H�U�H��H�E�H�E�H��HE�H�E��    H�u�H�E�H�E�����UH��H����H�����I��     L�H��     H�H�U�H�p0     H�H�R H�U�H�p0     H�H�U�H��H�P H�E�H� H��tH�E�H� H�P�H�E�H������UH��H����H�����I��     L�H�p0     H�H�R H�U�H�p0     H�H�U�H��H�P �����UH��AWH��(��H�����I��     Lډ}�H��     H�    H���������H�<I�׸    H�u�������H�������UH��H�� ��H�����I�D     L�H�}�u�H��     H�H�E��}� u,H�E�H���������H��H��H�E�H���H�E�H� H��u�����UH��H����H�����I��     L؉}��u��U��    ����UH��AWSH����H�����I��     L۾   �   I��H���������H��ЉE�}��u"H���������H�<I��H��������H����NH���������H�<I�߸    H�u�������H��ҋE��ЋE������M����Ɖ�H�"�������H���H��[A_]���UH��AWH����H�����I��     L�H��0     H�H�JH��0     H�H��0     H�H��t H��0     H�H�J�H��0     H�I��H�o@������H��ҐH��A_]���UH��H����H�����I�E     L؉}��4 �    �u�E���6   �C   �E��@   �E������@   �����UH��H����H�����I��     Lى}��H��0     H�    H��0     H�    H� �������H�H��������H�H�P�}� t"�6   �C   �d   H���������H�����2   �C   �����UH��H����H�����I�E     L�H�}�H��0     H�U�H���H��0     H�H��u됐����UH��H����H�����I��     L؉}��E�'  �}� u/�怃}� xZ�d   ���E��E�����uH�E��P��U���u��9�}�u3�怃}� x(�d   ���E��E�����t�E��P��U���u����������UH��H����H�����I�Q     L؉}��   H��������H��ЋE��d   �����UH��H����H�����I�	     Lؿ    H��������H��и`   ���E��E�����UH��SH����H�����I��     L��E�d   �    H���������H��҈E���    H���������H��҈E�}� x�}��t�E�P��U��u����H��[]���UH��AWSH����H�����I�:     Lۉ��E�   I��H��������H��и�   �d   �   I��H��������H����E�`   �H��[A_]���UH��AWH����H�����I��     Lؿ    I��H��������H��Ҹ`   ���E��E�H��A_]���UH��SH����H�����I�o     L۸    H�0�������H��҈E�}�u�    �$�}��u��������   H���������H����H��[]���UH��SH����H�����I��     L�H��0     ��PH��0     �����   ���=  ��t
��t(�/  �`   ���E��E��H��0     ��)  H��0     �������t(�`   ���E��E� �����H��0     ���   �`   ���E��E�H��0     ���   H��0     ����� ��t%�`   ���E��E� �����H��0     ���`   ���E��E�H��0     �H��0     ���xH��0     �����@��u�    H���������H���H��0     �    ��`   ���E�H��0     �    ��H��[]���UH��AWS��H�����I�F     L�H��0     H��H��0     �H��0     H�ʉH��0     H��HH��0     �H��0     H�)щʉPH��0     H�H��0     H��R�PH��0     �H��0     H��҉PH��0     H�� ��yH��0     H��     �HH��0     H�� ��H��������H��@9�v!H��������H��PH��0     H��H��0     H��@��yH��0     H��@    �JH��0     H��@��H��������H��@9�v"H��������H��PH��0     H��PH��0     H��PH��0     H�� �։�I��H��������H���H��0     H�H��0     H��   H��H��I��H�o�������H��А[A_]���UH��AWSH����H�����I�
     L�H��0     �    H��0     �    H��0     � H��0     �   H��0     �   �   I��H�R�������H���H��0     H�H��0     H��   �    H��I��H��������H��п   I��H�R�������H���H��H�0�������H�H�H�0�������H�H� H��H��0     H�H��0     H��   �    H��I��H��������H���H��������H��@���H��0     H��H��������H��@���H��0     H��PH��������H��PH��0     H���PH��0     H�H��������H��R�PH� �������H�H���������H�H�P`�   I��H��������H��и    �d   �    I��H��������H��и`   ���E��E�E�M��   I��H��������H��и`   �d   �   I��H��������H����E�`   �   I��H��������H��и�   �d   �    I��H��������H��п�   H���������H���I�߸    H�5�������H��ҿ�   H���������H���I�߸    H�5�������H��ҿ�   H���������H���I�߸    H�5�������H��ҿ�   H���������H���I�߸    H�5�������H��ҿ�   H���������H���I�߸    H�5�������H��ҿ   H���������H���I�߸    H�5�������H��ҿ�   H���������H���I�߸    H�5�������H��ҿ�   H���������H���I�߸    H�5�������H��ҐH��[A_]���UH��AWH����H�����I��     Lؿ    I��H��������H��Ҹ`   ���E��E�H��A_]���UH��AWH����H�����I��     L؉��U�   I��H��������H����E�`   �H��A_]���UH��SH����H�����I�I     L۸    H��������H��҈E�}�u�    �$�}��u��������   H�U�������H����H��[]���UH��AWSH����H�����I��     L۸`   ���E��E�E�}�;u8H�(�������H�H�H���������H�H�H��     �    ��  �E��y�}�t�}�uFH��     �    �3�}�*t�}�6u'H��     �   H��     �    �  �E��x�}�EuO�}��u3H��     ��PH��     �H��     �    �L  H��     �    �6  H��     ���tH��     ���u+�E�H��������H�H����H��0     ��  H��     ����a  H��     �    �E��P��   ��P�`  ��M�(  ��M�N  ��Ht��K��  �;  H���������H�H� H�ƿ   I��H���������H���H���������H�H� H�ƿ[   I��H���������H���H���������H�H� H�ƿA   I��H���������H����  H���������H�H� H�ƿ   I��H���������H���H���������H�H� H�ƿ[   I��H���������H���H���������H�H� H�ƿB   I��H���������H����/  H���������H�H� H�ƿ   I��H���������H���H���������H�H� H�ƿ[   I��H���������H���H���������H�H� H�ƿC   I��H���������H����   H���������H�H� H�ƿ   I��H���������H���H���������H�H� H�ƿ[   I��H���������H���H���������H�H� H�ƿD   I��H���������H����&�E�H��������H�H����H��0     �H��0     ���t9H���������H�H�H��0     ���H�։�I��H���������H���H��0     � H��[A_]���UH����H�����I�^      L�H��0     � H��     �    H��     �    H��     �    H��     �    �H� �������H�H��������H�H�B�]���UH��AWSH����H�����I���     L�H�}�H�h�������H�H��0     H��   I��H�R�������H���H��0     H�H��0     H�H��I��H��d������H���H��H��0     H�H�E�H��0     H�H��0     H�H��H�f������H��АH��[A_]���UH��H����H�����I���     L�H�}�H�E��@����H�E��P�H�E��@% @  ��u�H�E��@�����H�E��P�H�E��@% �  ��u�����UH��H����H�����I�s�     L�H�}��H�E��@% �  ��u�H�E��@����H�E��PH�E��@����H�E��P�����UH��AWSH����H�����I��     L�H�}�H�u�H�E�H��H�������H���H��0     H���H�E�H�E��@    H�E� ���   �    H��I��H��������H���H�E� ��   H�E�PH�E��@    H�E�@���   �    H��I��H��������H���H��0     H�H��   H��0     H�H�E�H��H��������H��АH��[A_]���UH��H��H��H�����I���     L؉}�H�uЉ׉�D��L�M��UD�E@�}�@�u�f�M�f�U�D�U��E�    H�U�H�U�H�U�H��@H�U�H�U��'H�U��J����JH�U��J�ᏈJ�U؉у�H�U������J��	�JH�U��B H�U��M̈JH�U��M��JH�P�������H��M�Hc�H��H�H�� ���t����   �  �Eȉ�H�E��PH�E���H�E��PH�E�H����H�E��PH�E�H����H�E��PH�E��@@H�E�H����H�E��PH�E�H�� ��H�E��P	H�E�H��(��H�E��P
�E�f����H�E��P�E���H�E��P�E�f����H�E��P��   �Uȉ�H�U��J�U�f����H�U��JH�P�������H��U�Hc�H��H�H��� �E��E���H�E��P�E�����H�E��PH�E��@@H�E�� �H�E��@ H�E�H����H�E�PH�E�H����H�E�PH�E�H����H�E�PH�E���H�E�PH�E��@ H�E��@ H�E��@ �E���H�E�P	H�E��@
 H�E��@ ������UH��H����H�����I�`�     L�H�}�H�u��U�H�E���H�E����   H�E�ǀ�       H�E�ǀ�       �E�%��? ��H�E��с���? ���   ��  ��	ʉ��   H�E����   f��?�f���   H�E����   �ʀ���   �����UH��H��(��H�����I���     L�H�}��u�H�U��D�ϋu�M�U�D�U���U���U܉ʈU��U��у�H�U�΃��
���	�
H�P�������H��U�Hc�H��H�H�� � ����H�E����������	ʈ�E����H�E���������	ʈ�E�����H�E�������	ʈ�E܃���H�E�у��P���	ʈP�E؃���H�E����P���	ʈPH�E��P����PH�E��P����PH�E��P���P�E ��H�E�f�PH�E�U(�PH�E��@��   H�E�PH�E��@    �����UH��AWSH��@��H�����I�$�     L�H�}ȉ�H�M���UĈE��E�    �E�    H�E��@����H�Eȋ ��H�E�H�U�H�E�j jj j A�    A�    �   �    H��H�G������H���H�� H�E��@��H�E�H�E��@����H�H��	����H�Eؾ    H��I��H��������H���H��0     H�H�Eغ�  H��H��H��������H���H�E�H�E�H�E�� '�E�����H�EЉу��P���	ʈPH�E��P�ʀ�PH�E��@��U�H�EЈP�E�   ����Љ�H�EȉP8�AH�Eȋ@ ����t/H�h�������H�<I�߸    H�u�������H��Ҹ�����  �E�H�Eȋ@ %�   ��t	�}�?B ~��}�@B u/H���������H�<I�߸    H�u�������H��Ҹ�����   H�EȋP8�E�   �����!Ѕ�t<H�Eȋ@%   @��t�H���������H�<I�߸    H�u�������H��Ҹ�����g�H�E��@=   t,H���������H�<I�߸    H�u�������H��Ҹ�����,H��0     H�H�E��@����H�E�H��H����    H�e�[A_]���UH��AWSH��0��H�����I�X�     L�H�}ȉu�H�Eȋ@(�E�E������E�E���E��E�    �E�    �E�    �}�t
������R  �}�t
������B  H�Eȋ@$=  ��  �E�   �E�   H�E�H��0     H��    �����H��H��������H��ЋE�H�P�������H��M�Hc�H��H�H�� �H��0     ���   ��%   ��t�0   ��   H�P�������H��U�Hc�H��H�H���HH��0     �Db��������H�P�������H��M�Hc�H��H�H���P�E�H�P�������H��M�Hc�H��H�H���H��0     �Dx��H�P�������H��M�Hc�H��HʉBH�P�������H��U�Hc�H��HЋ@H��0     �Tz�����H�P�������H��M�Hc�H��HȉP�  H�Eȋ@$=���   �E�   �E�   H�E�H��0     H��    �����H��H��������H��ЋE�H�P�������H��M�Hc�H��H�H�� ��E�H�P�������H��M�Hc�H��H�H���H�P�������H��U�Hc�H��H�H���@   H�P�������H��U�Hc�H��H�H���@0   H�P�������H��U�Hc�H��H��@    �~H�Eȋ@$=<�u�E�   �E�    �`H�Eȋ@$=i�u�E�   �E�    �B�E�    �E�    �Eĉ�H��������H�<I�߸    H�u�������H��Ҹ�����  H�(      �E�H�H�H�Eĉ�H��������H�<I�߸    H�u�������H��ыE�H�P�������H��M�Hc�H��H�H��0�BH�P�������H��U�Hc�H��H�H��0�@H�P�������H��M�Hc�H��H�H���B�E�H�P�������H��M�Hc�H��H�H��0�BH�P�������H��U�Hc�H��HЋ@   ���H�P�������H��M�Hc�H��HȉP�    H��0[A_]���UH��SH��(��H�����I���     L�H�}�H�E؋ �����E�U�H�P�������H��P�E�    �d�E�H�H��H��H��H�E�H�H�E�H��H��H��������H��ЋE�H�H��H��H��H�E�HE��H��H��
������H��ЃE��E�;E�|��    H��([]���UH��AWSH��@��H�����I���     Lۉ}�H�u�H�U��M�L�E�H�P�������H��U�Hc�H��HЋ@��x
�������  �E�    �E�    H�E��@����H�E�� ��H�E�H�U��u�H�E�j jj j A�    A�    �   H��H�G������H���H�� H�E��@��H�E�H�E��@����H�H��	����H�Eؾ    H��I��H��������H���H�P�������H��U�Hc�H��H�H��� �EȍP�H��0     H�H�E�H��H��H��������H���H�P�������H��U�Hc�H��H�H�� � ��t
��tu�   H�P�������H��U�Hc�H��H�H���@��u?�E���H�M�H�u؋E�j RI��A�    �%   �   ��H��������H���H���E������3  H�P�������H��U�Hc�H��H�H���@��u
������  �������   �E�   ����Љ�H�E��P8�H�E��@ ����t
�������   �E�H�E��@ %�   ��t	�}�?B ~ˁ}�@B u
������   H�E��P8�E�   �����!Ѕ�tH�E��@%   @��tո�����e�H�E��PH�P�������H��M�Hc�H��H�H��� �E�9�t�    �-H��0     H�H�E��@����H�E�H��H����H��    H�e�[A_]���UH��AWSH��@��H�����I���     Lۉ}�H�u�H�U��M�L�E�H�P�������H��U�Hc�H��HЋ@��x
�������  �E�    �E�    H�E��@����H�E�� ��H�E�H�U��u�H�E�j jj j A�    A�   �   H��H�G������H���H�� H�E��@��H�E�H�E��@����H�H��	����H�Eؾ    H��I��H��������H���H��0     H�H�P�������H��M�Hc�H��H�H����Uȉ���H�U�H��H����H�P�������H��U�Hc�H��H�H��� �EȍP�H��0     H�H�E�H��H��H��������H���H�P�������H��U�Hc�H��H�H�� � ��t
��tu�   H�P�������H��U�Hc�H��H�H���@��u?�E���H�M�H�u؋E�j RI��A�    �5   �   ��H��������H���H���E������  H�P�������H��U�Hc�H��H�H���@��u
�������   �������   �E�   ����Љ�H�E��P8�H�E��@ ����t
������   �E�H�E��@ %�   ��t	�}�?B ~ˁ}�@B u������oH�E��P8�E�   �����!Ѕ�tH�E��@%   @��tո�����=�H�E��PH�P�������H��M�Hc�H��H�H��� �E�9�t�    ��    H�e�[A_]���UH��SH��H��H�����I�<�     Lۉ}�H�u��U�H�M�H�E��E��E�    �E�    �E����E�H�E�H�E��E�    �   H�P�������H��U�Hc�H��H�H����E������E܋U�H�E�H�<�U�H��0     H��M�Hc�H��H��H�4�E�I���   ��H�3������H��ЉE�E�H�P�������H��U�Hc�H��H�H��� ��    �E�ЉE��}� t�E��n�E��E�9E��6����Eȃ��E؃}� tL�U�H�E�H�<�U�H��0     H��M�Hc�H��H��H�4�M؋E�I����H�3������H��ЉE�E�H��H[]���UH��SH��H��H�����I���     Lۉ}�H�u��U�H�M�H�E��E��E�    �E�    �E����E�H�E�H�E��E�    �   H�P�������H��U�Hc�H��H�H����E������E܋U�H�E�H�<�U�H��0     H��M�Hc�H��H��H�4�E�I���   ��H�h������H��ЉE�E�H�P�������H��U�Hc�H��H�H��� ��    �E�ЉE��}� t�E��n�E��E�9E��6����Eȃ��E؃}� tL�U�H�E�H�<�U�H��0     H��M�Hc�H��H��H�4�M؋E�I����H�h������H��ЉE�E�H��H[]���UH��H����H�����I��     Lى}�}���   H�P�������H��U�Hc�H��H�H�� �@�����E�H�P�������H��U�Hc�H��H�H�� �@�����E�H�P�������H��U�Hc�H��H�H�� �@�����E�H�P�������H��U�Hc�H��H�H�� �@�����E�������UH��H����H�����I�3�     L؉}�H�P�������H��U�Hc�H��H�H�� �@�����E��E�������UH��SH����H�����I���     Lۉ}��#�E��H��������H��Ѓ���t�   �#�E��H��������H���%�   ��u��    H��[]���UH��SH����H�����I�`�     Lۉ}��#�E��H��������H��Ѓ���t�   �#�E��H��������H���%�   ��t��    H��[]���UH��SH����H�����I���     Lۉ}��#�E��H��������H��Ѓ���t�   �!�E��H��������H��Ѓ���u��    H��[]���UH��SH����H�����I�t�     Lۉ}��#�E��H��������H��Ѓ���t�   �!�E��H��������H��Ѓ���t��    H��[]���UH��SH����H�����I���     Lۉ}�u��E��H�������H���H�P�������H��U�Hc�H��H�H�� �@�P�E��E��H��������H��АH��[]���UH��H����H�����I�z�     Lى}�H�P�������H��U�Hc�H��H�H�� �@���E��E��E��E�����H�P�������H��u�Hc�H��H�H�� �R��E�%�   H�P�������H��M�Hc�H��H�H�� �R�����UH��H����H�����I���     L؉}�H�u��U�H�P�������H��U�Hc�H��H�H�� �P�E����H�E�H����fm�����UH��H����H�����I�c�     L؉}�H�u��U�H�P�������H��U�Hc�H��H�H�� �P�E����H�E�H����fo�����UH��H����H�����I���     L؉}��u��U�M�D�E�D�M�U�H�P�������H��u�Hc�H��H�H��0�Q�U�H�P�������H��u�Hc�H��H�H���Q�U�H�P�������H��u�Hc�H��H�H�� �Q�U�H�P�������H��u�Hc�H��H�H�� �Q�U�H�P�������H��u�Hc�H��H�H�� �Q�UH�P�������H��M�Hc�H��H�H��0������UH��SH����H�����I���     Lۉ}�E��H�z������H��ЋE��H�������H���H�P�������H��U�Hc�H��H�H�� �@�P�    �H�P�������H��U�Hc�H��H�H�� �@�P�    �H�P�������H��U�Hc�H��H�H�� �@�P�    �H�P�������H��U�Hc�H��H�H�� �@�P�    �H�P�������H��U�Hc�H��H�H���@���H�P�������H��M�Hc�H��H�H�� �R���E��H��������H��ЋE��H�������H��ЋE��   ��H��������H��ЋE��H��������H����E�@B ��E��H��������H���%�   ��t�E�P��U��u����E��H��������H��ЉE��}� u
�    �   H�P�������H��U�Hc�H��H�H�� �@�����E��E�E�H�P�������H��U�Hc�H��H�H�� �@�����E��E�E�}�u�}��u�   �>�}�iu�}�u�   �+�}� u�}� u�   ��}�<u�}��u�   ��    H��[]���UH��AWSH����H�����I�$�     Lۉ}�H�u��E��H� ������H��Ѓ��w  ��H��    H�n� H�H�c� H�>���E��H�8�������H�<I�߸    H�u�������H���H�M��E�   H�Ή�H�,������H��ЋE��H�������H��ЋE��H�
������H���H�E�� f��y���  ��   H�P�������H��U�Hc�H��H�H�� �H�E�H�   � ��%   ��t�0   ��   H�P�������H��U�Hc�H��H�H���HH�P�������H��U�Hc�H��H�H���@    H�P�������H��U�Hc�H��H�H���    �  �E��H�I�������H�<I�߸    H�u�������H��ҋE쾡   ��H��������H��ЋE��H��������H��ЋE��H�������H���H�M��E�   H�Ή�H�,������H��ЋE��H�������H��ЋE��H�
������H���H�E�� f��y�   ����  H�P�������H��U�Hc�H��H�H�� �H�P�������H��U�Hc�H��H�H���@   H�P�������H��U�Hc�H��H�H���@    H�P�������H��U�Hc�H��H�H���    �   �E��H�\�������H�<I�߸    H�u�������H������E��H�m�������H�<I�߸    H�u�������H�����H�P�������H��U�Hc�H��H�H�� �     �E��H���������H�<I�߸    H�u�������H��Ґ�    H��[A_]���UH��AWSH����H�����I�S�     Lۉ}�u�H�U�H�P�������H��U�Hc�H��H�H���@��0�  ��0��  ����  ����  �E��H�P�������H��U�Hc�H��H�H�� �@�P���H�E���H�P�������H��U�Hc�H��H�H�� �@�P���H�E�H����H�P�������H��U�Hc�H��H�H�� �@�P���H�E�H����H�P�������H��U�Hc�H��H�H�� �@�P���H�P�������H��U�Hc�H��H�H���@����H�E�H������	Ѓ�@H�P�������H��M�Hc�H��H�H�� �R���H�P�������H��U�Hc�H��H�H���PH��2     �9���  H�P�������H��U�Hc�H��H�H�� �PH��2     �9��Q  �E��H��������H���H�P�������H��U�Hc�H��H�H���@H��2     �H�P�������H��U�Hc�H��H�H�� �@H��2     ���  H�P�������H��U�Hc�H��H�H�� �@�P�    �H�E�H����H�P�������H��U�Hc�H��H�H�� �@�P���H�E�H�� ��H�P�������H��U�Hc�H��H�H�� �@�P���H�E�H��(��H�P�������H��U�Hc�H��H�H�� �@�P���H�P�������H��U�Hc�H��H�H�� �@�P�E��H�E���H�P�������H��U�Hc�H��H�H�� �@�P���H�E�H����H�P�������H��U�Hc�H��H�H�� �@�P���H�E�H����H�P�������H��U�Hc�H��H�H�� �@�P���H�P�������H��U�Hc�H��H�H���@����@H�P�������H��M�Hc�H��H�H�� �R���H�P�������H��U�Hc�H��H�H���PH��2     �9���   H�P�������H��U�Hc�H��H�H�� �PH��2     �9���   �E��H��������H���H�P�������H��U�Hc�H��H�H���@H��2     �H�P�������H��U�Hc�H��H�H�� �@H��2     ��/�E��H���������H�<I�߸    H�u�������H���������H��[A_]���UH��SH��(��H�����I���     Lۉ}�u�H�U�H�M�H�P�������H��U�Hc�H��H�H�� � ����  ����  ��t
��t�|  ������w  H�U��M�E�Ή�H��&������H���H�P�������H��U�Hc�H��H�H���@��t���  �   H�P�������H��U�Hc�H��H�H���@��t��0t�7�E�    ��H��������H�����E�$   ��H��������H��А�E��H�������H��ЋE��H�������H��Ѕ�t
������   H�P�������H��U�Hc�H��H�H���H�M؋E�H�Ή�H�,������H��ЋE��H�������H��ЋE��H�
������H��Ѕ�t���������������������    H��([]���UH��SH��(��H�����I���     Lۉ}�u�H�U�H�M�H�P�������H��U�Hc�H��H�H�� � ����  ����  ��t
��t��  �������  H�U��M�E�Ή�H��&������H���H�P�������H��U�Hc�H��H�H���@��t���y  �  H�P�������H��U�Hc�H��H�H���@��t��0t�7�E�0   ��H��������H�����E�4   ��H��������H��А�E��H�������H��ЋE��H�������H��Ѕ�t
�������   H�P�������H��U�Hc�H��H�H���H�M؋E�H�Ή�H��������H���H�P�������H��U�Hc�H��H�H���@��t��0t�7�E��   ��H��������H�����E��   ��H��������H��А�E��H�������H��ЋE��H�
������H��Ѕ�t���������������������    H��([]���UH��AWSH�� ��H�����I���     Lۉ}܉u؉UԋUԋu؋Eܹ    ��I��H���������H��ЉE�H��     H��U�f��E�����H��     H�f�P�Uԋu؋Eܹ   ��I��H���������H��ЉE�E�����H��     H��P
�E�����H��     H��PH��     H��U�P	H��     H��@
<u,H��     H��@<uH�3     �   �  H��     H��@
<uNH��     H��@<u8H�3     �   H���������H�<I�߸    H�u�������H�����H��     H��@
<u)H��     H��@<uH�3     �   �qH��������H�<I�߸    H�u�������H���H�#�������H�<I�߸    H�u�������H���H�?�������H�<I�߸    H�u�������H������Uԋu؋Eܹ   ��I��H���������H��ЉE�E������Uԋu؋E�A�ȹ   ��I��H�P�������H���H��     H��@
<��   H��     H��@<��   �Uԋu؋Eܹ   ��I��H���������H��ЉE�E�% �  ��tR�Uԋu؋Eܹ   ��I��H���������H��ЉE�E�����Uԋu؋E�A�ȹ   ��I��H�P�������H���H��     H��@
<�C  H��     H��@<�)  �Uԋu؋Eܹ@   ��I��H���������H��ЉE�E� � ����Uԋu؋E�A�ȹ@   ��I��H�P�������H��ЋUԋu؋Eܹ   ��I��H���������H��ЉE�E�% �  ��tR�Uԋu؋Eܹ   ��I��H���������H��ЉE�E�����Uԋu؋E�A�ȹ   ��I��H�P�������H��ЋUԋu؋EܹH   ��I��H���������H��ЉE�E�����Uԋu؋E�A�ȹH   ��I��H�P�������H��ЋUԋu؋Eܹ<   ��I��H���������H��ЉE�H��     H��U�P/�E�����H��     H��P0�Uԋu؋Eܹ   ��I��H���������H��Љ�H��     H��P�Uԋu؋Eܹ   ��I��H���������H��Љ�H��     H��P�Uԋu؋Eܹ   ��I��H���������H��Љ�H��     H��P�Uԋu؋Eܹ   ��I��H���������H��Љ�H��     H��P�Uԋu؋Eܹ    ��I��H���������H��Љ�H��     H��P�Uԋu؋Eܹ$   ��I��H���������H��Љ�H��     H��P#�    H�� [A_]���UH��AWSH�� ��H�����I�L�     L�H�`�������H�<I�߸    H�u�������H��Һ   �    H�3     H�<I��H��������H��п   I��H�R�������H���H�E�   I��H�R�������H���H��     H��   I��H���������H��ЉE܃}��u'H���������H�<I�߸    H�u�������H������E��ЋE������M����Ɖ�H�]0������H��ЉE܃}� t'H���������H�<I�߸    H�u�������H�����H��     H��@�����H��     H��@��u��  ��    �H��     �H��     H��@�����H��     H��@��u��  ��    �H��     �H��     H��@�����H��     H��@��u�p  ��    �H�     �H��     H��@�����H��     H��@��u�v  ��    �H��     �H��     H��@�����H��     �H��     H��@#�����H�     �H�3     ���t���  �  H���������H�<I�߸    H�u�������H���H��     ���H��     ���H��     �H��RA��A���    �    �   �    I��H��������H���H��H��     ���H��     ���H��     �H��RA��A���    �   �   �   I��H��������H���H��H��     �����H��     ���H�     �H��RA��A���   �    �   �   I��H��������H���H��H��     �����H��     ���H�     �H��RA��A���   �   �   �   I��H��������H���H���E�    �"H�U��E�H�։�I��H��"������H��ЃE��}�~�H���������H�� ����H���������H��H�H�������H���   H���������H�<I�߸    H�u�������H���H�     ���H�Eй    �    H��I��H��S������H���H�E�H��I��H�0 ������H����'H��������H�<I�߸    H�u�������H������    H�e�[A_]���UH��AWSH��0��H�����I���     Lۉ}܉u�H�U�H�M�H�E�H�E�H�3     ���t
��t�   �E�    �gH�3     �E�H�H�H��H�H����E���H�E�H��E�Hc�H�E�HEܾ   ��I��H� ,������H��Ѕ�t������H�E��E�9E�w��5H�M��U�H�uЋE܉�I��H��������H��Ѕ�t��������������    H��0[A_]���UH��AWSH��0��H�����I���     Lۉ}܉u�H�U�H�M�H�E�H�E�H�3     ���t
��t�   �E�    �gH�3     �E�H�H�H��H�H����E���H�E�H��E�Hc�H�E�HEܾ   ��I��H��-������H��Ѕ�t������H�E��E�9E�w��5H�M��U�H�uЋE܉�I��H�K������H��Ѕ�t��������������    H��0[A_]���UH��H����H�����I���     Lظp   ���E��E��E��M���E��p   �����UH��H����H�����I�L�     Lظp   ���E��E��E��e��E��p   �����UH��H����H�����I��     Lظ
   �p   �q   ���E��E�%�   ����UH��AWSH����H�����I���     L�H�)�������H�<I�߸    H�u�������H��ҿ(   I��H�R�������H���H�;     H�H�;     H��(   �    H��I��H��������H���H�;     H��@$   H� �������H�H�o@������H�H�P@�    H�a>������H��Ҹ�   �p   �q   ���E��E�E踋   �p   �E��"�q   �    H��>������H��ҐH��[A_]���UH��SH����H�����I���     Lې�    H��>������H��҅�u�    �p   �q   ���E��E��P��H������������q   ���E��E����H�;     H���?��   �p   �q   ���E��E��P��H������������q   ���E��E���H�;     H���?�P�   �p   �q   ���E��E�P��H������������q   ���E��E���H�;     H����PH�;     H��HH�;     H��P$H�;     H�ʉPH�;     H��@��~H�;     H��@    �   �p   �q   ���E��E��H��     ��H��[]���UH��AWH����H�����I���     Lڸ    �怿
   I��H�������H�����H��A_]���UH��H����H�����I�V�     L؉}��U�U�H��;     H�H�H�E�H�E��U������UH��H����H�����I��     L؉}��f�U�U�H��;     H�H�H�E�H�E��U�f������UH��H����H�����I���     L؉}�u�U�H��;     H�H�H�E�H�E��U������UH��H����H�����I�d�     L؉}�U�H��;     H�H�H�E�H�E�� ����UH��H����H�����I��     L؉}�U�H��;     H�H�H�E�H�E�� ����UH��H����H�����I�Ի     L؉}�U�H��;     H�H�H�E�H�E�� ����UH��H�� ��H�����I���     L؉}�u�U�M�H��;     H�H�U�H�(;     ���H��    H�U�H��    H�(;     ���H��    H�U�Hʋ
�U����H�(;     ���H�<�    H�U�H�	�
H�(;     ���H��    H�U�Hʋ
�U����H�(;     ���H�<�    H�U�H�	�
H�(;     ���H��    H�U�Hʋ
�U����H�(;     ���H�<�    H�U�H�	�
H�(;     ���H��    H�U�HʋH�(;     ���H�4�    H�M�H�U��H�(;     ��JH�(;     ������UH��SH����H�����I��     L۾    �   H��B������H��и    H�OB������H��Ґ�   H��C������H���������u�  �   H��B������H��и    H�OB������H��Ґ�   H��C������H���������tᐐH��[]���UH��AWSH��P��H�����I��     L۾   �   I��H���������H��ЉE�H��;     �    H��;     �H�,;     �H�(;     �    H��;     �    H��;     �H��;     �H��;     �    H�<;     �    �}��u/H�@�������H�<I�߸    H�u�������H��Ҹ�����%  H���������H�<I�߸    H�u�������H��ҋE��ЋE������M����Ɖ�H�X������H��ЉEă}� t/H���������H�<I�߸    H�u�������H��Ҹ�����  H�8;     �   H�8;     �H�,;     ��׹    ��H��;     H�4I��H��S������H���H��;     H�H��H�0;     H�H�0;     H��@��H�0;     H��@����H� �������H�<I�߸    H�u�������H���H��;     H��   �    I��H��^������H���H��;     H��    �    H��I��H��������H���H��;     H�H��   H��;     H�H��;     H��    �    I��H��^������H���H��;     H��   �    H��I��H��������H��и    H�F������H��Ҿ    �    H�BC������H��о    �L   H��B������H��о    �\   H��B������H��о    �p   H�BC������H��о    �t   H�BC������H��о    �`   H�BC������H��о    �d   H�BC������H��о    �h   H��B������H��о    ��   H�BC������H��о   �   H�BC������H���H��;     H�H��I��H��d������H���H�E�H�E��ƿ  H�BC������H���H�E�H�� �ƿ  H�BC������H��о   �$  H��B������H���H�E�   H�E��ƿ�   H�BC������H���H�E�H�� �ƿ�   H�BC������H��о    �4   H�BC������H��о    �H   H��B������H��о    �L   H��B������H�����    H�OB������H��ҿL   H��C������H���������u̾    �\   H��B������H�����    H�OB������H��ҿ\   H��C������H���������u�H��;     H�H��I��H��d������H���H�E�H�E��ƿ@   H�BC������H���H�E�H�� �ƿD   H�BC������H���H��;     H�H��I��H��d������H���H�E�H�E��ƿP   H�BC������H���H�E�H�� �ƿT   H�BC������H����E�    �(�    �   �    �    H�gD������H��ЃE��}�	~Ҿ
   �H   H��B������H��о
   �Z   H��B������H��о �  �J   H��B������H�����    H�OB������H��ҿJ   H��C������H�����% �  = �  uǾ    �J   H��B������H�����    H�OB������H��ҿJ   H��C������H���f��xѾ �  �X   H��B������H��п\   H��C������H��Ѓ�������ƿ\   H��B������H��пL   H��C������H��Ѓ�������ƿL   H��B������H����*�J   H��C������H��и    H�OB������H��ҿX   H��C������H��Є�t�H�0;     H��@��H�0;     H��@��H�0;     H��@D��H�0;     H�D�@H�0;     H��@��H�0;     H��@��H�0;     H�� ��WV��H�8�������H�<I�߸    I�u�������I�A��H��H�0;     H��@N��H�0;     H��@M��H�0;     H��@L��H�0;     H��@J��H�0;     H��@H��A��A����H���������H�<I�߸    I�u�������I�A���E�    ��   �    H�H;     H�<I��H��������H��и    H�\Y������H���H�E�H���������H�<I�߸    H�u�������H��ҹ   �   �    �    H��Y������H��Ѕ�t%H���������H�<I�߸    H�u�������H���H�E�� ��H���������H�<I�߸    H�u�������H���H�E�� �����E�H�E�� ���E��E���H���������H�<I�߸    H�u�������H��ҋE��   �   �ƿ    H��Y������H��Ѕ�t%H���������H�<I�߸    H�u�������H���H�E�� ��H���������H�<I�߸    H�u�������H��ҋE��   �   �ƿ    H��Y������H��Ѕ�t%H���������H�<I�߸    H�u�������H���H�E�� �����E�H�E�� ���E��U��E���H���������H�<I�߸    H�u�������H����E�    �E�    �E�   ��  �EԹ	   �   �ƿ    H��Y������H��Ѕ�t%H���������H�<I�߸    H�u�������H��Ҹ    H�\Y������H���H�E��E�P�U�H�U��H�H;     H�Hى�H�E�� ����+  H�E�� ���  H�E�� ������uR�}� uL�E�   �E�H��;     ��EԉE��E���H��������H�<I�߸    H�u�������H����   H�E�� ������uS�}� uM�E�   �E�H��;     �H��;     ���H�'�������H�<I�߸    H�u�������H����XH�E�� ������uG�E�H�<;     �H�<;     ���H�=�������H�<I�߸    H�u�������H������E��U��E��9E��)����E��H�R�������H�<I�߸    H�u�������H����E�    �@H�H;     �E�H�Hڋ���H�f�������H�<I�߸    H�u�������H��҃E��E�;E�|��
   I��H���������H��ЋE���H�j�������H�<I�߸    H�u�������H��ҋE��    �  �ƿ    H��Y������H����E�    ��    H�OB������H��҃E��}�c~�E��    �  �ƿ    H��Y������H���H�E�� ��H��������H�<I�߸    H�u�������H��ҋE��   �   �ƿ    H��Y������H���H�E�� ��H���������H�<I�߸    H�u�������H���H�<;     ���   �
  �ƿ    H��Y������H���H�<;     ��    �
  �ƿ    H��Y������H���H�E�� ��H���������H�<I�߸    H�u�������H����E�    ��   �U��E�Љƿd   H��b������H��ЋU��E�й    �   �ƿ    H��Y������H���H�E�� ��H���������H�<I�߸    H�u�������H��ҋU��E�й   �   �ƿ    H��Y������H���H�E�� ��H���������H�<I�߸    H�u�������H��҃E��}��'����    H��`������H��ҋE���H�0^������H��и    H�e�[A_]���UH��AWSH�� ��H�����I��     Lۉ}܉u؉UԋUԋu؋Eܹ   ��I��H���������H��ЉE�E�����Uԋu؋E�A�ȹ   ��I��H�P�������H��ЋUԋu؋Eܹ   ��I��H���������H��ЉE�E�����H�,;     ��Uԋu؋Eܹ   ��I��H���������H��ЉE�H��;     �E��Uԋu؋EܹD   ��I��H���������H��ЉE�E� ���Uԋu؋E�A�ȹD   ��I��H�P�������H��и    H�� [A_]���UH��H����H�����I���     L�H��;     H�H��H�E�H�E�����UH��SH��(��H�����I�W�     Lۉ}܉u؉UԉM�H�(;     �    H��;     H�H�E�    �H   H��B������H��о    �L   H��B������H�����    H�OB������H��ҿL   H��C������H���������u̾    �Z   H��B������H��о    �\   H��B������H�����    H�OB������H��ҿ\   H��C������H���������u̹    �    �    �    H�gD������H��ЋMЋUԋu؋E܉�H�gD������H��й    �    �    �    H�gD������H��о   �H   H��B������H��о   �Z   H��B������H��о �  �J   H��B������H�����    H�OB������H��ҿJ   H��C������H�����% �  = �  uǾ    �J   H��B������H�����    H�OB������H��ҿJ   H��C������H���f��xѾ �  �X   H��B������H��п\   H��C������H��Ѓ�������ƿ\   H��B������H��пL   H��C������H��Ѓ�������ƿL   H��B������H����E�d   �>�J   H��C������H��и    H�OB������H��ҋE�P��U��u�������X   H��C������H��Є�t��    H��([]���UH��SH��(��H�����I��     Lۉ}܉u؉UԉM��E�    �E���	E�E���	E�E���	E�E�	E�   �h   H��B������H��ЋE�ƿ`   H�BC������H��о   �h   H��B������H����E�    �E�    �9�h   H��C������H���������t!�    H�OB������H��҃E��}�c~����}�d~������5�d   H� D������H��ЉE�   �h   H��B������H��ЋE�H��([]���UH��AWSH�� ��H�����I���     Lۉ}�H���������H�<I�߸    H�u�������H��ҋEܹ   �   �ƿ    H��Y������H��Ѕ�t*H���������H�<I�߸    H�u�������H�����  �    H�\Y������H���H�E�H��;     �@   H��;     �H�E� ��H� �������H�<I�߸    H�u�������H���H� �������H�<I�߸    H�u�������H��ҋEܹ   �  �ƿ    H��Y������H��Ѕ�t*H�?�������H�<I�߸    H�u�������H����  �    H�\Y������H���H�E�H�E� ��H���������H�<I�߸    H�u�������H���H�W�������H�<I�߸    H�u�������H���H��;     ��̰�E܉Ѻ   �ƿ    H��Y������H��Ѕ�t'H�c�������H�<I�߸    H�u�������H����F�    H�\Y������H���H�E�H�E� ��H���������H�<I�߸    H�u�������H��ҐH�� [A_]���UH��AWATSH��8��H�����I�*�     L�H��;     H�H�E�H�E�    H�E�H�E��E�   H�Eȉ�H�EЉH�E�H���     H�E�H�P�E��H�E�H���     �E��ƿ  H�BC������H��о C  �  H��B������H��о   �  H��B������H��о   �p   H�BC������H��о    �t   H�BC������H��о  �   H�BC������H��о   �4   H�BC������H����E�    ��    H�OB������H��҃E��}�c~�    H�OB������H��ҿt   H� D������H���A�Ŀp   H� D������H���D���H�{�������H�<I�߸    H�u�������H��ѐH��8[A\A_]���UH��H�� ��H�����I�R�     L؉}�u�H��;     �J   H��;     ��U��щU��U�Hc�Hi���QH�� ����)щʉU��M� �  �U��u�Ѻ   �    I��Y������J� �А����UH��H����H�����I���     Lظa   ���E��E����a   �����UH��H����H�����I�x�     Lظa   ���E��E�%�   �a   �����UH��H����H�����I�7�     L؉�f�E���   �C   ��E��B   ��E�f���B   �����UH��SH����H�����I��     Lۉ�f�E��E��H��c������H���H�=c������H��АH��[]���UH��AWSH�� ��H�����I���     L�H�}�H�E�H��@H�E�H�E�h   H��H�<     H�<I��H�o�������H���H�<     H�D(    H�<     �D8    H�<     �D<    H�<     �DH�<     �D@H�<     �DH�<     �DDH�<     �DP   H�<     �DT   H�<     �DX��� H�<     �D\    H�0�������H�H��H�<     H�T`�    H��h������H��ҐH�� [A_]���UH��H����H�����I�5�     L�H�}��u�U��U�H�<     �T�U�H�<     �TH�<     �TH�<     �TH�<     �D8    H�<     �D<    H�<     �TH�<     �T@H�<     �TH�<     �TDH�<     �DL    H�<     �TLH�<     �THH�<     H�U�H�T0�����UH��H����H�����I�)�     L�H�}�H�u��U�H�<     �T��H�U�H��H�U�H�H��    H�<     H�D0H�H�E������UH��H��0��H�����I���     L�H�}�H�u��U�H�M�H�U�H�U�H�<     �T��H9U�}KH�<     �T��H9U�}5H�<     �D��H�E�H��H�E�H�H��    H�E�HE܉������UH��AWH����H�����I��     L�H�<     H�T0H�U�H�<     H�T(H�U�H�<     �L@H�<     �TD��H�<     �L����H�u�H�M�H��I��H�o�������H��ѐH��A_]���UH��AWS��H�����I�s�     L�H�<     �T@H�<     �DD��H�<     �T����H�<     H�T0H�щ¾    H��I��H��������H���H�<     �DL    H�<     �DLH�<     �DH�[A_]���UH��SH��@��H�����I���     Lۉ}ԉuЉỦM�L�E�L�M�f�E�  H�E�H�@H�E؋EȉE�}�u�E�    �E�    �   f�E� H�E��@�ẺE��H�H� H�E�H�� f�E�H�E�� ���E��C�E�f#E�f��t.�UЋE��HcȋUԋE��H��U�H��H��H��f������H���f�e�m��}� y��E�H�E��@9E��i�����H��@[]���UH��SH����H�����I���     Lۉ}�}�
u9H�<     �DH    H�<     �DL�PH�<     �TL�E���  H�<     �DLH�<     �TT��H�<     �DD9�rH�<     �DL    H�<     �DHH�<     �TP��H�<     �D@9�r1H�<     �DH    H�<     �DL�PH�<     �TL�}���   H�<     �DH��t!H�<     �DH�P�H�<     �TH�PH�<     �DL��t>H�<     �DL�P�H�<     �TLH�<     �D@�P�H�<     �THH�X<     H�4H�<     H�D(I��H�<     �TXH�<     �DLH�<     �LT��A��H�<     �DHH�<     �LP���ǋE�I��щ�D��H�:i������H��Ѓ}�tH�<     �DH�PH�<     �TH�E�H��[]���UH��H��8��H�����I�Z�     L�H�}�H�uЉŰE����E�H�E�H�E�H�E�H�E��EH�E�� ��yH�E�� %��� ��H�E��H�E�H�E��H�U�H�BH�E�H�E�H�HH�M����E��P��U���u�H�E�����UH��AWSH�� ��H�����I���     L�H�}�H�E�H�  H�E�H�E�H��<     H��H��<     H�H�@H��u�H��<     H�H�PH��H�PH��<     H�H�E��4H�E�H� H9E�uH��<     H�H�@    ��   H�E�H�@H�E�H�}� u�H�E�    �    H��I��H��������H���H�E�H�U�H�H�E�H�@    H��<     H�H�PH��<     H�H��<     H��BdH��<     H�H�E��H�E�H�@H�E�H�E�H�@H��u�H�E�H�U�H�PH��<     H�H�@    H�� [A_]���UH��H����H�����I�)�     L�H�}�H��<     H�H�RH��u�H��<     H�H�JH��H�JH��<     H�H�U�H�U�H�U��   H�U�H�H9U�udH�U�H�RH��txH�U�H�JH�U�H�JH�U�H�B    H��<     H�H�U��H�U�H�RH�U�H�U�H�RH��u�H�U�H�M�H�J�!H�U�H�U�H�U�H�RH�U�H�}� �p�����H��<     H�H�@    �����UH��AWSH�Ā��H�����I��     L�H��x����H��<     H�H�@H��u�H��<     H�H�PH��H�PH��<     H�H�@H�x<     H��H  H�x<     H�H� H���  H�x<     H�H� H��H��<     H��H��<     H�� ��u�H��<     H�����H��<     H�H   H�E�H��x���H�E�H��<     H��@��H�E�H��<     H��@ ��H�E�H��<     H��PH��������H��@��H��<     H��@ �����H�E�H��<     H��@��H�E�H��<     H��@��H�E�H�E�H�E�H�U�H�E�H�H��������H��@��H9�~,H�U�H�E�H�H��������H��@��H)�H�E�H)�H�E�H��<     H��     H��������H��@��H9E�~%H�x<     H�H�@H�x<     H��y  �E�    �>  �E�H�H�U�H��H��H��H�E�H�H�E�H��������H��@��    �E���H�E�H�H�E�H�H�E�H�E؃�H��t0H�E�H��H�E�H�e�H�E؉�H�E�)ЉE��   +E�H�HE�H��<     H��@d��tU�E�Hc�H�E�H�H��������H��@��$��H9�}pH�E��    H�M�H�E�H��H��I��H���������H����CH��������H��P�E�9�v+H�E��    H�M�H�E�H��H��I��H���������H��ЃE��E�H�H9E������H�x<     H�H�@H�x<     H�H�x<     H�H�������H��<     H�H�@    �H��[A_]���UH��AWSH��0��H�����I���     L�H�}�H�u�H���������H��@4����  H��<     H�E�H�H�@�������H�H� �PH��<     H��PH�@�������H�H� �H��<     H��P H���������H�H�E��E�    �  �E�    ��   H��<     H��P�E��ЋE�Љ�H�E�H�� ���E܃}�uPH��<     H��P�E�Љ�H��<     H��P �E�Љ�H�E�H�������I��H�>g������H����T�}�uNH��<     H��P�E�Љ�H��<     H��P �E�Љ�H�E�H���  I��H�>g������H��ЃE�H��<     H��P�E�9������E�H��<     H��P�E�9��������H��0[A_]���UH��AWSH�� ��H�����I��     L�H�p<     �    �H��������H�H�@(H�¾   �    I��H��^������H���H�x<     H��   �    I��H��^������H���H�E�H�¾   �    I��H��^������H��и    ��H�x<     H��   �    H��I��H��������H���H�x<     H�H��<     H�H�`�������H��     H��������H�H�@0H�E�H��������H�H�@(H�E�H��������H��P@H��������H��@D��H��������H��@���E܋U�H�E�    H��I��H��������H���H�E��@   H�E��@   ����H���������H�H�H���������H��H��H��H��H��H�H�H��H)�H��u��H�E�H��H��o������H���H�U�H�E�H��H��H��s������H��АH�p<     ���u�H�p<     ��PH�p<     ��U�H�M�H�E�H��H��I��H���������H���H�p<     �    �'�����UH��AWSH��0��H�����I�p�     L�H�}�H�u�H�E�H�E��E�    H�E�   H���������H�4H��I��H�G�������H��Ѕ�u	�E�   �|H�E�   H���������H�4H��I��H�G�������H��Ѕ�u	�E�   �CH�E�   H���������H�4H��I��H�G�������H��Ѕ�u	�E�   �
�    �   �K  I��H�R�������H���H�E�H�EغK  �    H��I��H��������H���H�E��@    �    I��H�R�������H���H�U�H�BH�E�ǀ+      H�E��@"�U�H�E؉PH�E�H�@�    �    H��I��H��������H���H�E�H��0[A_]���UH��H����H�����I�ą     L؉}�H�u�H�U����H�U��R9�sH�U��J#H�U��R9�r"H�U��B'    H�U��J'H�U��J#H�U�f�  H�U��R��u&H��<     H��U�H�Ή�H�0z������H���H�E�H�PH�E��@#��H�H�E�H�PH�E�H�@�U��H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  �E�����UH��H�� ��H�����I���     L�H�}��E�    H�U�R����   H�U�R'�JH�U�J'��H�U�J#H�U�R'9�r�H�U�H�JH�U�R'��H��H�H�U�H�JH�U�H�R��҉U��}���   H��<     H��U�H�Ή�H�0z������H����   H�E�@��tH�E�@��uiH�E�@#��u������ZH�E�P'H�E�@#9�r������AH�E�H�PH�E�@'��H�H�E�H�PH�E�H�@� ���E�H�E�@'�PH�E�P'�E�����UH��H��0  ��H�����I�^�     L�H������H������H������H�E�H������H�E�H������H�E��E�    �?H�E�� ��u�E�Hc�H�E�H��  �H�E�H�PH�U��U�Hc�H�U�H�� ��E��}�_~��E�    �-H�E�H�PH�U��H�E�H�PH�U�� 8�t�   ��E��}�_~͸    ����UH��AWH����H�����I�x�     L�H�}�H�u�H�U��R��H�U����H�U�H��H��   I��I�5<������I�A��H��A_]���UH��AWSH��P��H�����I��     L�H�}�H�u�H�U��M�L�E�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H�R�������H���H�E�H�Eغ    �    H��I��H��������H��ЋU�H�E��@ H�M��	��H�M؉�I��H�5<������H��ЉE�}� t�E��   �E�    �7�E���Hc�H�E�H�H�E�H��H��H��|������H��ЉE�}� t�E��}�?~����}� u8�}�?2�E���Hc�H�E�H�H�EȺ�   H��H��I��H�o�������H���H�E�H��I��H���������H��ЋE�H��P[A_]���UH��AWSH��`��H�����I���     L�H�}�H�u�H�U��K  I��H�R�������H���H�E�H�EкK  �    H��I��H��������H���H�E��PH�E��@ ��H�EЉP�    I��H�R�������H���H�U�H�BH�E��PoH�EЉ�+  H�E��PH�EЉ�/  H�E��P H�EЉ�3  H�E��H�EЉ�?  �    I��H�R�������H���H�U�H��C  H�E�H��C  �    �    H��I��H��������H���H�E��@k�E�    I��H�R�������H���H�E��E������E�    �E�    ��  �   I��H�R�������H���H�U�H��C  �M�Hc�H��H�H�H�E�H��C  �U�Hc�H��H�H� H�E�H�E��   �    H��I��H��������H����E�    �>  H�E��@ �E��H�E��@�H�E��P�E�H�H�4�    H�E�H�ʉH�EЋ�;  �PH�EЉ�;  �E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E�;E�tu�E�H�U����H�U�H��H�¾   I��H�5<������H��ЉE��}� t:H�E�H��I��H���������H���H�E�H��H�V�������H��и    �   �E��E�H�E��@�����E�    ��U�E�H��    H�E�HЋ �E�}��u	�E�������E��}��  ������}��t�E��}��  ������H�E�H��I��H���������H���H�E�H��`[A_]���UH��AWSH��P��H�����I�}     L�H�}�H�u���   I��H�R�������H���H��<     H�H��<     H���   �    H��I��H��������H��п   I��H�R�������H���H�E�H�E�   �    H��I��H��������H���H�E��   �    H��I��H��������H����E�   H���������H�� ���E�H�U�H�E�H��H��H�z}������H��ЉE�}� tFH��<     H�H��I��H���������H���H�E�H��I��H���������H��и    ��   H��<     H�H�M�H�U�H�u�I�ȹ    H��H��}������H��ЉE�}� tCH��<     H�H��I��H���������H���H�E�H��I��H���������H��и    �pH��<     H�H�U�H�M�H��H��H�n������H���H�E�H��<     H�H��I��H���������H���H�E�H��I��H���������H���H�E�H��P[A_]���UH��AWSH�� ��H�����I��z     L�H�}�H�}� u
�������   H�E�H�@H��I��H���������H����E�    �TH�E�H��C  �U�Hc�H��H�H� H��t?H�E�H��C  �U�Hc�H��H�H� H��I��H���������H��ЃE��}��  ~���H�E�H��C  H��I��H���������H���H�E�H��I��H���������H��и    H�� [A_]���UH��AWH��(��L�����I��y     M�H�}؉u�H�E؋�;  �E�9�vH�}� u
������   H�E�H��C  �Eԍ��  ��H���
H�H��H�H� H�E�Eԙ���%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E؋�3  H�u؋�?  ����M��H�5<������L���H��(A_]���UH��AWSH�� ��H�����I��x     L�H�}�H�uпK  I��H�R�������H���H�E�H�E�K  �    H��I��H��������H���H�E��@    �    I��H�R�������H���H�U�H�BH�E�ǀ+      H�E��@"H�E��@   H�E�H�@�    �    H��I��H��������H���H�E�H�� [A_]���UH��H�� ��H�����I��w     L�H�}�H�u��E�    H�E�H�E��   H�E�� ��H�E��@9�sH�E��P#H�E��@9�rH�E��@#    H�E�f�   H�E�H�PH�E��@#��H�H�E�H�PH�E�H�PH�U�H�U�H�R� �H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  �E��}��E����E�����UH��H�� ��H�����I��v     L�H�}�H�u��E�    H�E�H�E�H�E��@'�PH�E��P'H�E��P'H�E��@9�rH�E��@'   �H�E��P#H�E��@'9�r�H�E��@'�P�H�E��P'�JH�E�H�PH�E��@'��H�H�E�H�PH�E�H�PH�E�H�HH�M���H�E��@'�PH�E��P'�E��}�~��E�����UH��H�� ��H�����I��u     L�H�}���U��E�E��E�H�E�H�E��H�E�H�PH�U��U��m��}� u�H�E�����UH��H��8��H�����I��u     L�H�}�H�uЉŰẺE�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M����E��P��U���u�H�E�����UH��H��0��H�����I�u     L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E��  H�E�����UH��H����H�����I��t     L�H�}�H�E�H�E��H�E�H�E�� ��u�H�E�H+E�����UH��H�� ��H�����I�Gt     L�H�}�H�u�H�E�H�E�H�E�H�E��3H�E��H�E�� 8�u!H�E�� ��H�E�� ��Ѕ�u�    �'H�E�H�PH�U��H�E�H�PH�U�� 8�t����������UH��H��(��H�����I��s     L�H�}�H�u��U��E�    �/�E�Hc�H�E�H���E�Hc�H�E�H�� 8�t�   ��E��E�;E�|ɸ    ����UH��H�� ��H�����I�7s     L�H�}�H�u�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E�����UH��AWSH��@  ��H�����I��r     L�H������H������H������H������H�E�f�E�  �E� �E�    ��  �E�Hc�H������H�� ����%��  �E��E�Hc�H������H�� ����X�� �.  ��H��    H��l H�H��l H�>��H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E��EӈE�H�U�H�E�H��H��H���������H���H�E��  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�U�H�E�H��H��H���������H���H�E��%  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E�H�������E�H�։�I��H�w�������H���H������H�E�H��H��H���������H���H�E��}  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E��E�H������H�։�I��H�w�������H���H������H�E�H��H��H���������H���H�E���   H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EԋE�H�������   H�Ή�I��H��������H���H������H�E�H��H��H���������H���H�E��*H�E�H���������H�4H��H���������H���H�E��9�E�Hc�H������H�� �E�H�U�H�E�H��H��H���������H���H�E萃E��E�Hc�H������H�� ���	���H�U�H������H)�H��H��@  [A_]���UH��AWH����H�����I�Un     L؉}�U��I��H�Dj������H���H��A_]���UH��AWSH�� ��H�����I�n     L�H�}�H�}� tT�E�    �)�E�Hc�H�E�H�� ����H���������H��ЃE�H�E�H��I��H�a�������H��ЋU�9�w���H�� [A_]���UH��AWSH���  ��H�����I�ym     L�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�H��0����   �    H��I��H��������H���ǅ���   ǅ���0   H�EH�� ���H��@���H��(���H�����H�����H��0���H��H��I��H�)�������H��Љ�<���H��0���H��H��������H��Ћ�<���H���  [A_]���UH��AWSH�� ��H�����I�Ol     L�H�}�H�u�H�E�� ��u
�    ��   H�Eк   H���������H�4H��I��H�G�������H��Ѕ�u&H�U�H�E�H��H��I��H��x������H���H�E��zH�Eк   H���������H�4H��I��H�G�������H��Ѕ�u&H�U�H�E�H��H��I��H�=�������H���H�E��$H�U�H�E�H��H��I��H��������H���H�E�H�E�H�� [A_]���UH��AWH����H�����I�/k     L�H�}�H�}� u������H�U�H��I��H�V�������H���H��A_]���UH��H����H�����I��j     L�H�}�H�}� t7H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@����H�E��P������UH��H����H�����I�oj     L�H�}�H�u��U�}�tZ�}�|�}� t�}�t�nH�E���H�E��P#H�E���H�E��P'�RH�E��@#H�U��H�E��P#H�E��@'H�U��H�E��P'�(H�E���+  H�U�)Љ�H�E��P#H�E��P#H�E��P'�H�E��@#H�U��J�    ��Љ�H�E�f��    ����UH��H����H�����I��i     L�H�}�H�}� u�    �	H�E��@#������UH��AWH����H�����I�Ni     L؉}�H�u�H�U��R��tH�U��R��tH�U��R��u H�M��U�H�Ή�I��H�0z������H�����    H��A_]���UH��AWH��(��H�����I��h     L�H�}�H�E؋@��tH�E؋@��tH�E؋@��u$H�E�H��I��H�A{������H��ЉE�E���   H�E؋P#H�E؋�+  9�r
�������   H�E؋@����uIH�E؋@����H�E؉PH�E؋@#H�U؋r�    ���E�U�H�E؉�H��I��H�_�������H���H�E�H�HH�E�� ����H�U�f�2H��H�H�E�H�PH�E�H�@� ���E�H�E�� ��H�E؋@9�rH�E؋@����H�E؉PH�E�f�   H�E؋@#�PH�E؉P#�E�H��(A_]���UH��SH��H��H�����I�^g     L�H�}ȉuĉU�H�M�H�}� u�    �u�E�    H�E�H�E��E�    �FH�E�H��H�"�������H��ЉE܃}��u�E�    �u��0H�E�H�PH�U��U܈�E��E��E��E�9E�r��E�    �u�H��H[]���UH��AWH��(��H�����I��f     L؉}܋U����U�U܁��  ��t�E��M�H�U��ο   I��H��^������H���H�E�H��(A_]���UH��AWH����H�����I�1f     L�H�}�H�U�H��I��H�qa������H��ҐH��A_]���UH��AWSH��0��H�����I��e     Lۉ}�H�u��Uȃ}� u#H�E�H�E�H�E�H�PH�U�� 0H�E��  �  �ẺE��E�Hc�H�E�H�H�E��1�E����E��m��}�	~�7   ��0   �U��H�m���H�E�H�E�H;E�wŋE�Hc�H�E�H��  H�E�H�E��E�    �8H�E�� <0uH�E��"H�U�H�E�H��H��I��H��������H�����E��E�;E�|�H�E�H�E�H�E�H��I��H�a�������H��ЉE�   +E��M�H�U�Hщ¾    H��I��H��������H���H��0[A_]���UH��H��0��H�����I�}d     L؉}�H�u�H�E�H�E��E܉E��E�    �}� y,H�E�H�PH�U�� -�}�   �u�E�����E���E��؉E�H�E�H�E�M�Hc�Hi�gfffH�� ��������)�����)��ʉЍH0H�E�H�PH�U�ʈ�E�Hc�Hi�gfffH�� ����)ЉE�}� u��}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��H��H��H�����I�6c     L�H�}�H�u��U�H�E�H�E��E��E�H�E�H�E�H�E�H�E�H�E���H��uH�E���H��tW�E�����H�E�H�U�H��H����H��E܃���t*�E܃�A��H�U�H�E�H��H��D���H��H��H�U�H�E�H�E���   H�E� @ @@@`��   ��   ��   ��   �   �   �E����E؃}� tX�E�    �BH�E�H�U��@  �`  ( (H(P (X0++J+R +Z0H�E�@H�E�@�E��E�9E�w���w�E܃�?��t*�E܃�?A��H�U�H�E�H��H��D���H��H��H�U�H�E�H�E���f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ~ � � � � � � � � ~             ~ � � � � � � � � ~                 l � � � � | 8                   8 | � | 8                   < < � � �   <                < ~ � � ~   <                      < <              � � � � � � � � � � � � � � � �           < f B B f <           � � � � � � � � � � � � � � � �        2 x � � � � x             < f f f f <  ~               ? 3 ? 0 0 0 0 p � �              c  c c c c g � � �               � < � < �             � � � � � � � � � � �               > � >                  < ~    ~ <                f f f f f f f   f f              � � � {                | � ` 8 l � � l 8  � |                       � � � �              < ~    ~ <  ~              < ~                           ~ <                      �                         0 ` � ` 0                         � � � �                       ( l � l (                      8 8 | | � �                   � � | | 8 8                                                 < < <                  f f f $                             l l � l l l � l l           | � � � |   � � |               � �   0 ` � �             8 l l 8 v � � � � v           0 0 0 `                             0 0 0 0 0 0               0         0                   f < � < f                         ~                                    0                     �                                                           0 ` � �             8 l � � � � � � l 8              8 x       ~             | �    0 ` � � �             | �   <    � |               < l � �                 � � � � �    � |             8 ` � � � � � � � |             � �     0 0 0 0             | � � � | � � � � |             | � � � ~     x                                                       0                  0 ` 0                      ~     ~                     ` 0      0 `             | � �                       | � � � � � � � |              8 l � � � � � � �             � f f f | f f f f �             < f � � � � � � f <             � l f f f f f f l �             � f b h x h ` b f �             � f b h x h ` ` ` �             < f � � � � � � f :             � � � � � � � � � �             <         <                   � � � x             � f f l x x l f f �             � ` ` ` ` ` ` b f �             � � � � � � � � � �             � � � � � � � � � �             | � � � � � � � � |             � f f f | ` ` ` ` �             | � � � � � � � � |           � f f f | l f f f �             | � � ` 8   � � |             ~ ~ Z       <             � � � � � � � � � |             � � � � � � � l 8              � � � � � � � � � l             � � l | 8 8 | l � �             f f f f <     <             � � �   0 ` � � �             < 0 0 0 0 0 0 0 0 <               � � � p 8                 <         <          8 l �                                                   �       0                                     x  | � � � v             � ` ` x l f f f f |                   | � � � � � |                < l � � � � v                   | � � � � � |              6 2 0 x 0 0 0 0 x                   v � � � � � |  � x       � ` ` l v f f f f �                 8      <                        f f <       � ` ` f l x x l f �             8         <                   � � � � � � �                   � f f f f f f                   | � � � � � |                   � f f f f f | ` ` �             v � � � � � |                � v f ` ` ` �                   | � ` 8  � |              0 0 � 0 0 0 0 6                    � � � � � � v                   � � � � � l 8                   � � � � � � l                   � l 8 8 8 l �                   � � � � � � ~   �             � �  0 ` � �                 p                                        p         p                       v �                        8 l � � � �           RUN: kernel --> x86_64
 Setup LGDT ...\\
 Setup LIDT ...\\
 Setup Paging ...\\
 Setup MM ...\\
 Setup SMP ...\\
 Setup PIT ...\\
 Setup RTC ...\\
 Setup I965 ...\\
    Sirius OS (Kernel mode: AMD64 or x86_64)
CPU: %s
 stdin stdout stderr   Setup drivers de interface ...\\
 Keyboard ...\\
 Mouse...\\
 ATA ...\\
 Done
 Initialize....
 A: r+b launcher.bin fopen error launcher.bin
    Divide error
 Debug exception
 NMI Interrupter
 Breakpoint
 Overflow
 BOUND Ranger exception
   Invalide opcode (Undefined opcode)
     Device not avaliable (Not Math coprocessor
)    Double Fault (Erro de codigo)
  Coprocessor segment overrun (reservado)
        Invalide TSS (Erro de codigo)
  Segment not present (Erro de codigo)
   Stack segment fault (Erro de codigo)
   General protetion (Erro de codigo)
 Page fault (Erro de codigo)
 Intel reserved do not use 15
  x87 FPU Floating-Point error (Math fault)
      Alignment check (Erro de codigo)
 Machine check
        SIND Floating-Point exception
 Virtualization exception
 Intel reserved do not use 21
 Intel reserved do not use 22
 Intel reserved do not use 23
 Intel reserved do not use 24
 Intel reserved do not use 25
 Intel reserved do not use 26
 Intel reserved do not use 27
 Intel reserved do not use 28
 Intel reserved do not use 29
 Intel reserved do not use 30
 Intel reserved do not use 31
      CR2 = 0x%x - %x, CR3 = 0x%x, CR4 = 0x%x
 PYSICAL: %x %x
 PID:%d
        r+b open error "%s"
    ���������{������(~������_���������������������������ACPI MADT (Multiple APIC Description Table) ... \\ 
 APIC ACPI MADT not found!
 Found %d cores, IOAPIC %x, LAPIC %x
Processor IDs:  %d 
BSP ID: %d 
Initialize APs... \\ 
aprunning %x
 
Local APIC AP1: ID = %x  %x    Memory Map error, size > 1GiB
  Memory Map error, size > %d bytes, (0x%d bytes)
 Alloc Frame error
 FIXME frame APIC_LVT_PERFORMANCE
 APIC_LVT_LINT0
 APIC_LVT_LINT1
 APIC_LVT_ERROR
 Default LVT n: %d
        .�������J�������t���������������Ƞ��������������������*�������F�������b�������{�����������������������Null IRQ n: %d
 Erro IRQ%d
 APIC Global enable 0x%x
 stdin stdout stderr pipe _ cole _ Syscall %x error
        ? This help cd Change current directory clear Clear screen copy Copy file or directory date Date del Delete file or directory dir List directory echo This --- exit Exit shell help info This System information mov Move file or directory new New file or directory reboot Reboot system rename Rename file or directory shutdown     Shutdown your computer locally or remotely time Time version Shell version 

~ $  %c %s: command not found
 ~ $  Function not implemented
      Sirius OS (Kernel mode: AMD64 or x86_64)
CPU: %s
 Commands:
 SSE hardware not supported
 SSE is available
      Unclassified Mass Storage Controller Network Controller Display Controller Multimedia Controller Memory Controller Bridge device        Simple Communication Controller Base System Peripheral Input Device Controller Docking Station Processor Serial Bus Controller Wireless Controller Intelligent I/O Controllers  Satellite Communication Controller Encryption Controller Signal Processing Controller Processing Accelerator Non-Essential Instrumentation Co-Processor Unassigned Class (Vendor specific) Non-VGA-Compatible devices VGA-Compatible Device SCSI bus controller IDE controller (ISA Compatibility mode-only controller) IDE controller (PCI native mode-only controller)        IDE controller (ISA Compatibility mode controller, supports both channels switched to PCI native mode)  IDE controller (PCI native mode controller, supports both channels switched to ISA compatibility mode)  IDE controller (ISA Compatibility mode-only controller, supports bus mastering) IDE controller (PCI native mode-only controller, supports bus mastering )       IDE controller (ISA Compatibility mode controller, supports both channels switched to PCI native mode, supports bus mastering ) IDE controller (PCI native mode controller, supports both channels switched to ISA compatibility mode, supports bus mastering ) Floppy disk controller IPI bus controller RAID bus controller ATA Controller (Single DMA) ATA Controller (Chained DMA)  Serial ATA controller (vendor specific interface)       Serial ATA controller (AHCI 1.0 interface)      Serial ATA controller (Serial Storage Bus) Serial Attached SCSI (SAS)   Serial Attached SCSI (Serial Storage Bus)       Non-Volatile Memory Controlle (NVMHCI)  Non-Volatile Memory Controlle (NVM Express) Other mass storage controller Ethernet controller Token ring controller FDDI controller ATM controller ISDN controller WorldFip Controller PICMG 2.14 Multi Computing Infiniband Controller Fabric Controller Other Network controller      VGA Compatible controller (VGA Controller)      VGA Compatible controller (8514-Compatible Controller ) XGA controller  3D controller (Not VGA-Compatible) Other Display controller Multimedia video controller Multimedia audio controller (AC'97) Computer telephony device   Audio Device (Intel High Definition Audio (HDA) Controller) Other Multimedia controller RAM controller FLASH controller Other Memory controller Host bridge ISA bridge EISA bridge MCA bridge   PCI-to-PCI Bridge (Normal Decode)       PCI-to-PCI Bridge (Subtractive Decode) PCMCIA bridge NuBus bridge CardBus bridge        RACEway bridge (Transparent Mode)       RACEway bridge (Endpoint Mode)  PCI-to-PCI Bridge (Semi-Transparent, Primary bus towards host CPU)      PCI-to-PCI Bridge (Semi-Transparent, Secondary bus towards host CPU) InfiniBand to PCI host bridge Other Bridge Serial controller (8250-Compatible (Generic XT))        Serial controller (16450-Compatible )   Serial controller (16550-Compatible )   Serial controller (16650-Compatible )   Serial controller (16750-Compatible)    Serial controller (16850-Compatible)    Serial controller (16950-Compatible)    Parallel Controller (Standard Parallel Port)    Parallel Controller (Bi-Directional Parallel Port)      Parallel Controller (ECP 1.X Compliant Parallel Port)   Parallel Controller (IEEE 1284 Controller)      Parallel Controller (IEEE 1284 Target Device) Multiport Serial Controller Modem (Generic Modem) Modem (Hayes 16450-Compatible Interface)        Modem (Hayes 16550-Compatible Interface)        Modem (Hayes 16650-Compatible Interface)        Modem (Hayes 16750-Compatible Interface)        GPIB (IEEE 488.1/2) Controller Smart Card       Other Simple Communication controller PIC (Generic 8259-Compatible) PIC (ISA-Compatible) PIC (EISA-Compatible)  PIC (I/O APIC Interrupt Controller)     PIC (I/O(x) APIC Interrupt Controller)  DMA controller (Generic 8237-Compatible)        DMA controller (ISA-Compatible) DMA controller (EISA-Compatible)        Timer (Generic 8254-Compatible) Timer (ISA-Compatible) Timer (EISA-Compatible) Timer (HPET) RTC (Generic RTC) RTC (ISA-Compatible) PCI Hot-plug controller SD Host controller IOMMU     Other System peripheral controller Keyboard controller Digitizer Pen Mouse controller Scanner controller Gameport controller (Generic)  Gameport controller (Extended) Other input controller Generic Docking Station Other type of docking station 386 486 Pentium Alpha Power PC MIPS Co-processor    FireWire (IEEE 1394) controller (Generic)       FireWire (IEEE 1394) controller (OHCI) ACCESS Bus SSA USB (UHCI Controller) USB1.1 (OHCI Controller) USB2.0 (EHCI Controller) USB3.0 (XHCI Controller) USB Controller (Unspecified )    USB Device (Not a host controller) Fiber Channel SMBus InfiniBand IPMI Interface (SMIC) IPMI Interface (Keyboard Controller Style)      IPMI Interface (Block Transfer) SERCOS Interface (IEC 61491 CANbus iRDA controller Consumer IR controller RF controller Bluetooth Controller Broadband Controller       Ethernet Controller (802.1a – 5 GHz)  Ethernet Controller (802.1b 2.4 GHz)    Other type of wireless controller I2O Satellite TV controller Satellite audio controller Satellite voice controller Satellite data  controller  Network and Computing Encrpytion/Decryption     Entertainment Encryption/Decryption Other Encryption/Decryption DPIO module Performance counters Communication synchronizer Signal Processing Management        Other Signal Processing Controller Null PCI Listing devices:
 %s , B%d:D%d:F%d
 Other PCI Device ClassCode (%X), B%d:D%d:F%d
   panic: PCI Display Controller not found!
 Display Controller
   Graphic Native Intel, not found, device id %x, vendor id %x
    Checksum failed
 ACPI version 2.0,  ACPI version 1.0,  OEM_ID "%s"
 ACPI_Setup ... \\ 
 FACP acpi error
 DSDT _S5_ DSDT nao encontrado
 Use the 8042 keyboard controller to pulse the CPU's RESET pin
 HPET_Setup ... \\ 
      PCI PANIC: LPC Controller not found!
 LPC found
 Default Unknown IntelliMouse    1234567890-=	qwertyuiop[]
 asdfghjkl;'` \zxcvbnm,./                                                                                                                                                                                                           !@#$%^&*()_+	QWERTYUIOP{}
 ASDFGHJKL:"~ |ZXCVBNM<>?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          SATA SATAPI SEMB PM                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             sata(x) Read disk CMD ATA IDENTIFY error
 port(x) is hung 
     sata(x) read disk CMD ATA IDENTIFY error
       sata(x) read disk CMD ATA IDENTIFY error ---
 sata%d device not found
 sata%d device type: %s
  Uinidade%d PATA
 Uinidade%d PATAPI
 Uinidade%d SATA
 Uinidade%d SATAPI
 Uinidade%d Not found
   �0�������-������P0�������.������|0������PANIC,ATA Modo CHS not suport Unidade%d
        panic: RAID Controller
 IDE Controller not found!
 RAID Controller not found!
 AHCI Controller not found!
      Initializing the ATA Controller:
       PIC: Massa Storage Controller not found!
       PANIC: IDE/AHCI PCI Configuration Space
 IDE Controller:
 AHCI Controller:
     IDE or AHCI controller not found RTC install...\\
      PCI PANIC: Intel High Definition Audio (HDA) Controller not found!
     PCI Intel High Definition Audio Controller initialize
  PCI PANIC: Intel High Definition Audio (HDA) Controller error!
 Intel High Definition Audio Controller version %d.%d
   
GCAP:%x OUTPAY:%x INPAY:%x GCTL:%x WAKEEN:%x STATESTS %x GSTATUS:%x    
CORBWP:%x CORBRP:%x CORBCTRL:%x CORBSTATUS:%x CORBSIZE:%x
 Root Node:  error:
 %x
 Start Node %d, Parametro 5:   AFG: %d %d
 CORB/RIRB error:
 Output stream node %d
 Input stream node %d
 Beep Widget node %d
 
Numero de AFG: %d
 %x  HDA OUTPUT NODE: %d
 : %x
    Detalhes do amplificador de saida: %x
 Beep: %x
 : VOLUME %x
 HDA set output node
      CORB error: Get amplifier info
 Get amplifier info: %x, %d
     Set stream: stream 1 chanel 1
 CORB error: Set stream
 Set volume
 CORB error: Set volume
 %x %x
 stdin stdout stderr   %%      ��������\�������\�������\�������\�������\�������\�������\�������\�������\�������\�������P�������a�������\�������\�������\�������\�������a�������\�������\�������\�������\�������\�������\�������\�������\�������\�������ۓ������\�������	�������\�������\���������������std pipe                                                                                                                                                                                        Y%@     hE     �E     �+@     00E     �&E     �&@     n)@     �%@     %-@     5&@     �%@     -@     C-@     0E     �E     �+@     ,%@     80E     ��B     ��@     �,@     �E     0E     D&@     pE     �&@     xE     �-@      �A     0$E     })@     �&@     �+@     &&@     -@     @0E     �&@     J%@     H"E     �,@     &@     �%@     xE     �E     ,@     x"E     ;%@     �,@     �,@     %@     �#E     -@     p-@     �/E     g'@     H0E     ��A     a-@     �"E     �&E     �&E     �,@     �E     q&@     �%@     �A     �+@     �-@      $E     �+@     �#E     4-@     �%@     P0E     �,@     �#E     |E     �A     S&@     �%@     �-@     �E     �%@      E     E     X0E     `E     �-@     w%@     �,@     @$E     }iA     �)@     �)@     �%@     q,@     %@     h%@     �)@     �%@     �E      E     �%@     �-@     &@     �%@     �&@     �.E     R-@     �+@     b&@      �A     �,@     �,@                                              �A     .�A     ?�A     P�A     \�A     f�A     ��A     ��A     طA     ��A     (�A     H�A     p�A     ��A     ��A     ٸA     ��A     (�A     J�A     `�A     �A     ��A     ��A     չA     �A     �A     /�A     M�A     k�A     ��A     ��A     źA     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     ��@     !�@     y�@     Ѥ@     F�@     ǥ@     �@     ��@     �@     ^�@                      �A     �@     �A     �A     �@     �A     (�A     ��@     .�A     ;�A     O�@     @�A     W�A     �@     \�A     a�A     ��@     e�A     ~�A     &�@     ��A     ��A     ò@     ��A     ��A     `�@     ��A     ��A     �@     �A     ��A     �@     ��A     ѾA     ��@     վA     �A     K�@     �A     �A     �@     �A     �A     ��@     "�A     ;�A     4�@     H�A     s�A     ѭ@     x�A     }�A     n�@     ��A                     H�A     U�A     m�A     ��A     ��A     ��A     ��A     ��A     ��A     �A     �A     /�A     9�A     O�A     c�A     ��A     ��A     ��A     ��A     ��A                                                                                                                                                                                                                                                                                                                                                                     �A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �A         ;�A        V�A        l�A       ��A      ��A     
 ��A      X�A     � ��A     � �A     � `�A     � ��A       `�A       w�A       ��A       ��A     0 ��A       ��A      �A      @�A       k�A      ��A      ��A      ��A      � �A        *�A       >�A       T�A       d�A       s�A       ��A       ��A       ��A       ��A      � ��A        ��A       (�A       `�A       p�A      � ��A        ��A       ��A       ��A       �A      � D�A        `�A       o�A      � ��A        ��A       ��A       ��A       ��A       ��A      ��A       �A       %�A       2�A       H�A      p�A     @	 ��A     �	 ��A      
 �A      � ;�A        H�A       ��A       ��A       ��A       ��A        �A       H�A       p�A      ��A      ��A      �A     � @�A       n�A       ��A      ��A      ��A       �A      0�A       `�A       �A      � ��A        ��A       ��A       ��A        �A        (�A       P�A      ��A      ��A       ��A      ��A      ��A      �A       $�A      6�A       K�A       c�A       v�A      � ��A       	 ��A      	 ��A      	 ��A      	 ��A      	 ��A     	 �A      �	 '�A       
 >�A      �
 V�A        t�A       x�A       |�A       ��A        ��A      0 ��A      @ ��A        ��A       ��A       ��A       
�A       �A      $�A       =�A     0 V�A     � o�A     � ��A       ��A       ��A       ��A       ��A      ��A      �A       8�A      	 T�A        [�A       k�A       ��A       ��A       ��A        ��A      ! ��A      � �A        2�A        6�A       N�A       i�A       ��A        ��A       ��A      � ��A        �A       �A       1�A        L�A      � p�A         ��A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ��A     ��A     ��A     ��A                              �A     �A     �A     �A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    zR x�  ,      ����J	   E�CJ��4	�B�A�          L   ����B    E�Cy�     l   �����   E�C��,   �   �����   E�CC����B�A�          �   e���3    E�Cj�  $   �   x���s    E�CC��d�B�A�     ����   E�C	�$   $  �����    E�CC����B�A�   L  ���h    E�C_�    l  ����l    E�Cc� (   �  I���I   E�CC��:�B�A�       �  f����   E�CG��          �  �����    E�CF���A�       �����   E�CG��      ,   $  ����T   E�CI���=�B�B�A�      T   ��9    E�Cp�     t   ���    E�CI���   �  � ��G    E�C~�     �  � ��G    E�C~�     �  ��Z    E�CQ�    �  Y��2    E�Ci�       k��2    E�Ci�     4  }��,    E�Cc�     T  ���.    E�Ce�     t  ����    E�C�� (   �  ���   E�CG����B�A�   (   �  ���[   E�CG��H�B�A�   $   �  ����    E�CG����B�A�      [���    E�CF���A�   8  /	���    E�C�� (   X  �	���   E�CG����B�A�      �  d��~    E�Cu� (   �  ����   E�CG����B�A�   $   �  5��W   E�CE�H�A�       �  d���   E�C��          ��n    E�CE�_�A�    @  \���    E�CE���A�    d  ��K    E�CE�|�A�     �  6��i    E�CE�Z�A�   �  {��K    E�CB�    �  ���n    E�Ce� (   �  ���B   E�CG��/�B�A�   (     
���   E�CC����B�A�       D  ���\    E�CF�L�A�$   h  ����    E�CG����B�A�(   �  K���   E�CC����B�A�       �  � ��S    E�CF�C�A�    �  !��k    E�CF�[�A�     V!��=    E�Ct�  (   $  s!���   E�CG��r�B�A�      P  �#��F    E�C}�     p  �#��_    E�CV�    �  1$���    E�C��    �  �$��b    E�CY�    �  �$��@    E�Cw�     �  %��J    E�CA�      6%���    E�C��    0  �%���    E�C�� $   P  P&���   E�CE���A�       x  �(���    E�CE�{�� $   �  Z)���    E�CG����B�A�$   �  �)��k    E�CF�[�A�    ,   �  0*��<   E�CI���%�B�B�A�   ,   	  <-��(   E�CI����B�B�A�   (   L	  42���   E�CG����B�A�      x	  �5���   E�C��   �	  >���   E�Cw�    �	  kC��p    E�Cg�     (   �	  �C��   E�CJ���
�B�A�   (   
  �N��   E�CJ���B�A�       4
  ~Y��k    E�CF�[�A�    X
  �Y��X    E�CF�H�A�    |
  �Y��X    E�CF�H�A�   �
  -Z��u    E�Cl� $   �
  �Z���    E�CG��n�B�A�    �
  �Z��X    E�CF�H�A�$     [��|    E�CG��i�B�A�$   4  c[��|    E�CG��i�B�A�(   \  �[��G   E�CG��4�B�A�   $   �  �\���    E�CG����B�A�    �  x]���    E�CF���� $   �  �]��g    E�CF�W�A�       �  �^���   E�CJ��        Na��c    E�CF�S�A�    @  �a��c    E�CF�S�A�    d  �a��Z    E�CF�J�A�    �  b��c    E�CF�S�A�    �  Ab��Z    E�CF�J�A�    �  wb��c    E�CF�S�A�    �  �b��c    E�CF�S�A�$     �b���    E�CJ����B�A�(   @  �c��q   E�CG��^�B�A�       l  �d��c    E�CF�S�A�    �  /e��c    E�CF�S�A�    �  ne��c    E�CF�S�A�    �  �e��c    E�CF�S�A�    �  �e��c    E�CF�S�A�       +f��c    E�CF�S�A�    D  jf��Z    E�CF�J�A�    h  �f��c    E�CF�S�A�$   �  �f���    E�CG����B�A�,   �  cg���   E�CG��w�B�A�          �  �j��0    E�Cg�       �j��4    E�Ck�     $  �j��.    E�Ce�     D  �j��/    E�Cf�     d  �j��/    E�Cf�  $   �  k���    E�CG����B�A�   �  �k��|    E�Cs�    �  l��|    E�Cs�    �  tl��|    E�Cs�      �l��|    E�Cs� (   ,  ,m��   E�CG����B�A�      X  o���    E�C��    x  �o���    E�C��    �  �p���    E�C��    �  tq��   E�C�   �  cr��1    E�Ch�     �  tr��:    E�Cq�        �r��@    E�Cw�      (   <  �r���   E�CG����B�A�   (   h  -t���   E�CG���B�A�      �  �u���   E�C��   �  Qx��}    E�Ct�    �  �x��}    E�Ct�    �  y��    E�Cv�      jy��    E�Cv�    4  �y��    E�Cv�    T  (z��    E�Cv�    t  �z��+    E�Cb�     �  �z��?    E�Cv�     �  �z���    E�C��    �  Y{��+    E�Cb�     �  d{��?    E�Cv�       �{��F    E�C}�  $   4  �{���   E�CE���A�      \  }��1    E�Ch�     |  )}���    E�C��     �  �}��   E�CE���A�    �  �~��y    E�Cp�        �  0��P    E�CG� (     `���   E�CG����B�A�      0  ���T    E�CK�     P  M����    E�CE���A�(   t  �����   E�CG��w�B�A�      �  ]����    E�C�� (   �  	����   E�CG��}�B�A�      �  m����    E�C}�      Ӈ���    E�CF�       ,  n���j    E�Ca�    L  �����    E�C~�    l  ���W    E�CN�    �  V���b    E�CF�    �  ����r    E�Ci�        �  ���4    E�Ck�  $   �  �����    E�CG����B�A�      �����    E�CF���A�   8  ���^    E�CU�    X  I����    E�C��     x  ˋ��U    E�CL�        �  �����    E�C��    �  {���H    E�C�     �  ����J    E�CA� $   �  ͌���    E�CE�s�A�    $   $  '���y    E�CG��f�B�A�    L  x���T    E�CF�D�A�    p  ����u    E�CE�f�A�$   �  �����   E�CE���A�   (   �  ����'   E�CC���B�A�   (   �  ����+   E�CG���B�A�         ����T    E�CF�D�A�    8  ����U    E�CF�E�A�    \  ���u    E�CE�f�A�(   �  3���{   E�CG��h�B�A�      �  �����    E�C�� $   �  �����    E�CG����B�A�   �  ����t    E�Ck�      ���b    E�CY� (   4  C���   E�CG���B�A�      `  /����   E�C��   �  �����    E�C��    �  ;����   E�C}�(   �  �����   E�CG����B�A�   (   �  A����   E�CG����B�A�         ����    E�CE���A�(   <  ����5   E�CG��"�B�A�   (   h  ����O   E�CG��<�B�A�   $   �  �����   E�CE���A�   $   �  #����   E�CE���A�      �  �����    E�C��      Q���[    E�CR�     $  ����w    E�CE�h�A�    H  ߳��w    E�CE�h�A�    l  2���u    E�CE�f�A�    �  ����u    E�CE�f�A�    �  Դ���    E�CE�w�A�   �  6����    E�C��    �  ȵ��e    E�C\�      ���e    E�C\�    8  R���   E�C�$   X  J����   E�CE���A�   (   �  ����   E�CG����B�A�   (   �  ����b   E�CG��O�B�A�   $   �  �����   E�CE���A�   (      ����a   E�CE�R�A�       (   ,  ����H   E�CG��5�B�A�   (   X  �����   E�CG��}�B�A�   (   �  E���   E�CG���B�A�   (   �  /���   E�CG���B�A�      �  ���G    E�C~�     �  @���G    E�C~�       g���E    E�C|�  (   <  ����;   E�CG��(�B�A�   (   h  �����   E�CE���A�           �  O���O    E�CF��A�    �  z���Q    E�CH�    �  ����S    E�CJ�    �  ����N    E�CE�      ���H    E�C�     8  4���H    E�C�     X  \���G    E�C~�     x  �����   E�C��    �  
����    E�CE���A�(   �  ����2   E�CG���B�A�   (   �  ����P   E�CG��=�B�A�         ����@    E�Cw�  $   4   ����R   E�CE�C�A�   $   \   &���B   E�CE�3�A�   (   �   @����   E�CG����B�A�   ,   �   �����   E�CI�����B�B�A�       �   V����    E�C��        !  ����?    E�Cv�     $!  ����A    E�Cx�     D!  ���P    E�CG� $   d!  =���Y    E�CE�J�A�    (   �!  n���Y   E�CG��F�B�A�      �!  ����   E�C�   �!  ����s    E�Cj�    �!  �����    E�C��     "  Y����    E�CF���A�$   <"  �����    E�CC����B�A�    d"  j���
   E�CE���A�(   �"  P���V   E�CE�G�A�          �"  z����    E�C�� (   �"  �����   E�CG��|�B�A�       #  _���%   E�C�(    #  d ��   E�CG����B�A�   (   L#  <���   E�CG����B�A�       x#  ���   E�CG��      (   �#  y���   E�CG����B�A�      �#  �	��   E�C�    �#  �
��R   E�CI�       $  ���    E�C��     ,$  ���i    E�CF�Y�A�(   P$  '���   E�CG��x�B�A�   (   |$  ����   E�CG��n�B�A�   (   �$  ���g   E�CG��T�B�A�   $   �$  ��	   E�CG����B�A�$   �$  ����    E�CF���A�    $   $%  ����    E�CG����B�A�   L%  q��    E�C��    l%  Q���    E�C��    �%  ��b    E�CY�    �%  W��w    E�Cn�    �%  ���{    E�Cr�    �%  	��L    E�CC�    &  5���    E�C��    ,&  ���v    E�Cm�    L&  ��l    E�Cc� ,   l&  Q��t   E�CJ��^�B�A�           �&  ���H    E�CF�x�A� $   �&  ����    E�CG��}�B�A�(   �&  !��-   E�CJ���B�A�   (   '  " ��!   E�CG���B�A�       @'  !��Y    E�CF�I�A�   d'  L!��i    E�C`�    �'  �!���    E�C��    �'  S"��A    E�Cx�      �'  t"��~    E�CF�n�A�$   �'  �"��s   E�CF�c�A�       (  $���    E�CE���A�    4(  �$��o    E�CF�_�A�    X(  �$��L    E�CF�|�A� (   |(  %%��j   E�CG��W�B�A�       �(  c&��G   E�C>�       �(  �'���   E�C��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        GCC: (Ubuntu 9.3.0-17ubuntu1~20.04) 9.3.0                                      @                    �A                    �B                   ��B                   ��B                    C                    @E                                       ��                     ��  @                 �����            �     @                    =@             #      �@             0    ��                7      ��A             <      ��A             A      ʵA             F      ܵA             K      �A             P       �A             U      �A             Z      "�A             _      3�A             d      H�A             i      z�A             o      ��A             u      ��A             {      ��A             �      ��A             �      ¶A             �      ζA             �      ٶA             �      ߶A             �      �A             �      �A             �      ��A             �      �A             &   ��                �    ��                �     `@     �      �    ��                �    ��                �     � @           �    ��                     ��  @                 �����            �      �$@             �      �&@             �      '@                  {(@                  _)@                  �)@                  �*@                  �+@             )     ,@             1   ��                =     �A             C     �A             I     !�A             O   ��                V   ��                7      0�A             <      4�A             _   ��                7      ��A             <      ��A             A      ��A             F      лA             K      �A             P      �A             U      �A             Z      )�A             _      8�A             d   ��                l   ��                u   ��                7      X�A             <      x�A             A      ��A             F      ��A             z   ��                �   ��                �   ��                7      ȼA             <      ޼A             A      �A             F      ��A             K      �A             �   ��                7      ��A             <      ��A             �   ��                7      ��A             �   ��                �   ��                7      ŽA             <      ˽A             A      ҽA             F      ٽA             �   ��                7      ޽A             �   ��                7      �A             �   ��                     ��  @                 �����            �     @�@             �   ��                �     ��A             �     ��A             �     ��A             �     ��A             �     ��A                  ؿA                  
�A                ��                   ��                7      �A             <      1�A                ��                      ��A             '     ��A             .     ��A             5     ��A             <   ��                7      ��A             <      �A             A      0�A             C   ��                L   ��                S    �@     P       i    h�@     �      s    M�@     T       �    �@     �       7      p�A             <      ��A             A      ��A             F      ��A             K      ��A             P      ��A             Z      ��A             U      ��A             _      ��A             d      ��A             i      ��A             �   ��                �    @E            �    ��@     j       �    �@     �       �    ��@     W       7      7�A             �   ��                �    ��@     4       7      P�A             <      v�A             �   ��                �    ��@     �       �   ��                    ��@     J          ��                    G�@     '      !   ��                ,    DE            2    HE            <    LE            B    PE            H   ��                O     �A      �      Z    �A     �       o    ��@     t       x    �@     b       �    {�@           �    ��@     �      �    ,�@     �       �    ��@     �      �    e�@     �      �    1�@     �      �    �A     5      �     A     O      K       �B             P      *�B             U      @�B             Z      p�B             _      ��B             d      ��B             �   ��                �    �A     �          6A     b      7      ��B             <      ��B             A      ��B             F      �B             K      �B             P      X�B             &   ��                0    �#A     H      7      ��B             <      ��B             A      ��B             F      ��B             K      ��B             P       �B             U      P�B             Z      y�B             _      ��B             d      ��B             L   ��                R    �2A     E       i    `E            7      ��B             u   ��                {    �KA     P      7      ��B             <       �B             A      X�B             F      ��B             K      ��B             P      �B             U      T�B             Z      `�B             _      h�B             d      l�B             i      ��B             o      ��B             u      ��B             {      ��B             �      ��B             �      ��B             �      ��B             �      �B             �      �B             �       �B             �      G�B             �      Q�B             �      ^�B             �     x�B             �     ��B             �     ��B             �     ��B             �     ��B             �     ��B             �     �B             �   ��                �   ��                �   ��                �    2`A     �       �   ��                �   ��                7      �B             <       �B             A      '�B             �   ��                �   ��                   ��                   ��                    U�A     l       7      0�B             #   ��                7      @�B             <      D�B             +   ��                4   ��                     ��                A    ��B             W    5�A     H       _    Y%@             e    :VA     �       p    iC@     G       w    ~~A     {       ~    ��@            �    f�@     /       �    �@     c       �    ��@     �           hE            �    ��@     �      �    �2A     ;      �    �zA     �       �    0�@           �    ]TA     �      �    �E     
       �    �+@                  �A     -      �    00E            �    ��A     t          2�@     �           y�@     X       '    �7A     �      :    )A     e       H    �l@     @       ]    �Q@     ~       d    �.E            q    ��@     c       y    �&E            �    ($E            �    ��@     c       �    �m@     �       �     k@     F       �    �@             �    ,$E            �    ��@     �       �    WA     A       �    H�@     r            A     �           �&@                 ��@     �      "    n)@             '    �%@             -    w[@     K       3    !E            =    `$E            E    1�@     +       Q    \�@           ^    ��@     �      l    w�@     �      x    %-@             ~    XE            �    5&@             �    �%@             �    L$E            �    ("E            �    �@             �    -@             �    h$E            �    �C     8       �    �.E            �    C-@             �    0E            �    �E            �    wA     �       �    �"@     �           �+@                 ��A                 ,%@             &    80E            .     m@     J       D    �yA     �       T    ��B     �       e    �@     �       n    0E            t    )@     �      �    (E            �    ��@             �    �#E            �    �,@             �    �E     0       �    0E            �    ��@     U           ~A     w       �    ��B     �      �    D&@             �    ��@     �      �    pE            �    �7A     G       �    0"E            �    E            �    �&@             	    �a@     \       	    E            	    ��@           �	    }�A     �       %	    p�@     :       6	    A     u       C	    O�@     y       O	    ��@     �       Y	    8"E            e	    �E@     �      v	    ��@     �      �	    xE            �	    �-@             �	    �#E            �	    �A     o       �	    $E            c     �A             �	    0$E            �	    `0E            �     �E            �	    })@             �	    @E            �	    �K@     �           �!A     a      �    �r@     k       �	    ��B            �    	U@     W      �	    !�@     X       
    �g@     S       
    �&@             
    i�@     �       +
    ��@     }       6
    ^�@     �       C
    �+@             p	    OG@     [      J
    lE            S
    pE            \
    �A     G      a
    66A     Q       j
    &&@             p
    @"E            �     0E            {
    \A     �       �
    QD@     2       �
    �.E            �
     !E            �
    ��@     +       �
    % @     3       �
    ��@            �
    �9A     �       �
    -@             4    '�@     p       �
    @0E            �
    �&@                 J%@                 �@     u           d�@     |       ,    WYA           7     @E             @    	�@     }       L    �#E            U    �A           e    ��B     P       v    H"E            �    ��@     k       �    	�@     .       �    ѭ@     c       �    �`A     �      �    �,@             �    �.E            �    ��@     0       �    �ZA     �       �    �.E            �    �cA           �    x�@     1       �    @#E             �    P"E                ��@     �           �gA     �      '    &@             -    X"E            9    +A     w       G    ��@     {      X    \B@     9       ]    �@             O    �#E            e    �A     w       w    �%@             }    �k@     �       �    `X@     �      �    xE            �    YA     [       �    `"E            �    ƪ@     �      �    �E     h       �    �6@     �      �    A�@     �       �    �@     |       �    �h@     �           h"E                  E               (b@     �           չ@     4       %    (7A     H       -    4�@     Z       :    �q@     �       G    p"E            U    ,@             \    x"E            l    �"E            {    ;%@             �    �,@             �    l�@     |       �    �E            �    �@     |       �    cbA     %      �    �LA     @       �    �,@             �    {qA     �      �    K�@     c       M    ��@     �       �     pE             �    �M@     �      	    %@                 `#E                8$E                ��B            /    �A     �       c    �#@     h       5    �#E            :    -@             @    ��@     �       K    p-@             Q    �"E            \    �"E            i    n�@     c       u    ��@     Z       3    �/E     h           UWA     P       �    g'@             �    (0E            �    ��@     �       �
    H0E            �    @     B       �    ��A            �    �A     e       �    a-@             �    �"E            D     C             �    �&E            �     @             �     pE                 V�A     �      W    �&E                ��@     �           �.E     �       %    &�@     c       -    �D@     2       =    �Z@     �       S    �"E            _    �,@             d    �6A     N       (    `!E     �       m    �A             z    �E            �    �"E            �    �@     q          �0A           �    �\A     
      �    �"E            �    q&@             �    �C@     G       �    cZA     s       �    �PA     B      �    �"E            �    �%@             �    ��@     T       �    sA     �      E     C             g    �5@     �           �]A     V      �    `/E                �b@     �          ]�@     �       !    �"E            ,    �A             6    �-@     I      I    �A     v       �    �A     �      P    O�@     c       Y    �+@             `    �E            i    �E            r    �xA     	      }    �{A            �    �-@             �    E@     �       �    p$E            �    -�A     �       �     $E            �    �D@     ,       �    �"E            �    �+@             �    �@             �    �#E     8       ~    �vA     g      �    4-@             �    ,�@     �           �%@                 h/E                ��@           "    +�@     �      *    "4@     �      :    p/E            F    �E            I    :�A     !      V     �A             O    �}A     b       V    ;�@     H       c    �@     J	      h    �@             p    <$E            x    ��A     A       ~    �VA     ?       �    �5A     O       �    ��B            �    ǥ@     X       �    P0E            �    $E            �    �A     �       �    ^h@     =       �    �,@             �    [�A     Y       �     "E                4A     �          �A     �      "    �"E            -    \v@     (      ;    �nA     R      D    �#E            I    �@     Z       T     �A             [    Ѥ@     u       (    |E            l    2Z@     n       y    �A             �    S&@             �    �%@             �    (!E            �    &_@     �      �    +\@     K       �    EA     �       �    �-@             �    ��@     T       �     `E            �    �E            �    �"E            �    �%@             �     E            �    �"E            �    ��@     �      �    n�@     +          ��@     y       #    �"E            /    �{@     �      C     C             I    ��@     b       T    �@            b    7$@     l       l    ��A     s      r    E            x    �@     G      �    0!E            '    X0E            �    �QA     �      �    O
A     �      �    x/E            �    kM@     �       �    `E     
       �    �-@             �    p7A     H       �    N$E            �    �C@     Z       �    w%@                 fk@     _           �,@                 ��A                @     �      $    �n@     �      U     �A             ;    u[A     �       �    @$E            H    sL@     �       T    G�@     ^       g    <�A     ~       m    }iA     �      |    ��@     c       L    jR@     �      �    `�@     c       �    qq@     �       �    �)@             �    $E            �    ��@     @       �    m@             �    G�@     U       �    v\@     n       �    �)@             �    �D@     .       �    �%@             �    ��A     j      �    �\@     B          ��@     �           @2A     G            �@     c       '    �B@     �       2    2�@     �       C    <@     T      M    r:A     2      W    q,@             \    7�@     /       �     pE             e    %@             k    =*A     �      z    lA     �      �    �mA           �    ��A     i       �    ש@     g       �    ��@     |       �    �WA     Y      �    C@             *     @             �    �"E            �    h%@             �    �)@             �    �%@             �    �E            �    �#E            �    �|A     �       �    �@     �          H$E                ?�@     1            ^�@     �       /    �"E            ;    ò@     c       D    F�@     �       X     E            b    8!E            m     #E            y    ^l@     b       �    �1A     G       �    #E            �    �%@             �    #E            �    �g@     k       �    x$E            �    #E            �    �-@             �    eA     �      �    &@             �    0#E            �    �@                �%@                 f@                 �&@             !    �~A     L       (     @             /    �6A     S       8    +pA     �       E    �.E            )     @             K    �E            T    �E            ]    qA     i       n    �#E            w    �C             �    R-@             �    o�@     �       �    �+@             �    �#E            �    �[@     i       �    \�@     ?       �    *�@     ?       n     $E            �    �/E            �    @!E            �    X @     s           b&@                 �$E                ��A            (     s@     <      5     #E            A    �WA     Y       N    ��@           [    B�@     u       m    �/E            |    �/E            �    �@     |       �    �A     u       �     �A     h      �    4MA     R      �    ��@     F       �    �,@             �    �,@             �    �/A           �    Y�A     L       �    (#E            �    �/E            �    Jm@     �        setup.asm KERNELSTACK APsSTACK L1 copymem.loop main.c .LC0 .LC1 .LC2 .LC3 .LC4 .LC5 .LC6 .LC7 .LC8 .LC9 .LC10 .LC11 .LC12 .LC13 .LC14 .LC15 .LC16 .LC17 .LC18 .LC19 .LC20 .LC21 .LC22 gdt.c set_gdt tss.c idt.c set_gate_idt vetor.asm isr_jmp lvt_jmp lvt_jmp2 lvt0.loop iv timer1.loop __no_mult_task irq_jmp exception.c .LC32 .LC33 .LC34 data.c server.c mp.c delay.c paging.c mm.c cpuid.c msr.c lvt.c irq.c apic.c sleep.c thread.c exectve.c syscall.c asyscall.asm syscall_jmp console.c .LC35 .LC36 .LC37 .LC38 .LC39 .LC40 .LC41 exit.c sse.c pci.c .LC179 .LC180 .LC181 .LC182 i965.c cursor.c acpi.c acpi_set_virtual_addr init_rsdp acpi_check_header acip_init hpet.c timer_tick hpet_freq hpet_handler0 hpet_handler1 lpc.c lpc_pci_configuration_space pit.c pit_handler ps2.c kbdc_read mouse.c mouse_refresh keyboard.c shift caps_lock scaps count ahci.c _zhba_base sata_port_initialize stop_cmd start_cmd sata_port_confg sata_set_cfis sata_set_prdt sata_set_cmdHeader ahci_ata_indentify sata_identify ahci_read ahci_write ide.c detect_devtype set_ata_device_and_sector storage.c ata_pci_configuration_space rtc.c get_update_in_progress status.1539 hda.c hda_pci_configuration_space .LC23 .LC24 .LC25 .LC26 .LC27 .LC28 .LC29 speaker.c gui.c screen.c trans_memcpy font8x16.c std.c cfs.c pipe.c string.c vsprintf.c _vsputs_r stdio.c stdlib.c sse_memcpy.c _GLOBAL_OFFSET_TABLE_ putchar isr05 hda_volume mdelay strcpy enable_pipe fpu_restore cmd_date kbdc_wait gmbus_read rtc_setup pipe_open_file pci_scan_bcc_scc_prog hda_play_sound gdtr timer7 vsprintf keyboard_install syscall_window corb_write_command ata_pio_write read_ioapic_register v_pool corb_pointer cmd_mov ata_record_channel mouse_x cmd_del ioapic_umasked apic_initial_count_timer EnableSSE count_mouse DrawMouse turn_speaker_off hpet_sleep ata_soft_reset isr27 task_switch2 lvt1 isr13 cpuid alloc_pte dmavirt gmbus_reset pci_get_info mouse_handler acpi_enable irq12 ata_pci isr22 isr15 key_buffer context_rcx DisableSSE irq10 dmaphy ahci_type HDBARL irq14 screan_spin_lock thread_id ata_wait idt_install timer2 ascii_minusculas isr02 _stderr write_ioapic_register file_read_block fnvetors_handler cmd_info paint gdt_install call_loader int114 fadt irq8 server_id gid keyboard_write cmd_table isr23 setup_i965 kernelmouse hda_inl context_r12 pae_pde isr29 default_irq pae_pte exectve_child pci_check_vendor ata_wait_drq mouse_write setup_sse context_rax initialize_mm_mp setup_acpi dv_uid irq23 acpi_physical_init malloc eticks mouse2 fs_directory lvt2 mouse_position ram_setup exception_mensagem syscall_puts getapicbase isr31 disable_legacy_vga_emul enable_dac pci_scan_bcc timer6 ATA_BAR1 ATA_BAR4 itoa hda_outb isr21 context_ds clears_creen load_pae_page_directory_pointer_table hda_base alloc_pde disable_dpll load_ltr enable_plane hda_reset irq11 _stdin isr28 isr04 MOUSE_BAT_TEST pci_read_config_dword update_gui eh_frame disable_dac SLP_TYPa ata_bus_install fnvetors_syscall current_thread default_syscall sse_cw cmd_time window_add irq5 HDA_MEM_SIZE fpu_cw put_pixel_buff beep_node paint_desktop gmbus_write fb current_thread2 pit_enable paint_cursor isr20 context_rsi ata_wait_busy keyboard_handler done copymem ata_wait_not_busy isr14 apic_timer_umasked get_phy_addr user ata_status_read context_r9 console tss server pci_scan_class write_pci_config_addr setup_apic context_rdx core irq_function sse_cr hda_inb cmd_shutdown setup_ioapic context_rflag timer8 current_thread1 context_fxsave isr03 irq6 read_pci_config_addr CPUID_REQUEST syscall_readsector window_foco hda_response irq1 read_directory_entry cmd_new alloc_pages_setup isr01 mode first_time pci_class_names fseek xsdt irq18 acpi_probe irq17 context_cs context_rsp0 cmd_version cmd_clear set_speaker_frequence lvt0 paint_ready_queue setup_lpc font8x16 ata_pio_read irq16 thread_ready_queue ata_record_dev _start __end sse_memcpy kbdc_wait_ack hda_widget cmd_dir load_pml4_table cpuid_processor_brand context_cr3 irq9 hda_outl SavedFloats2 launcher context_rsp cmd_help draw_char_transparent context_fs isr26 udelay put_pixel hda_ic_verbe context_rbp isr11 mouse_read open_file_r glyph irq_install poweroff context_r8 _ap_stack exceptions_install memcmp cmd_copy timer5 ATA_BAR0 ATA_BAR3 file_close pipe_write irq19 page_install HBA_BASE fread timer_ticks enable_pae context_r15 timer4 RestoreSSE gtt irq13 syscall_function_handler isr12 HDA_STREAM_MEMORY exectve timings fault_exception RIRB_MEMORY no fopen memset kbdc_set_cmd main SaveSSE buttons ftell turn_speaker_on hda_wait pci_classes syscall_free_pages _stdout hpet_register ata_cmd_write apic_eoi_register irq2 fclose ioapic_base rtc_handler sata_write_sector context_ss create_thread std_getc rsdt cmd_reboot __data syscall_kbd_foco cpuid_vendor SavedFloats isr24 isr16 RAM_BITMAP lvt_install getmsr strcmp irq20 keyboard_read syspwd next_pid isr08 pml4e context_gs i965_pci_init mouse_install update_graphic_cursor context_r11 create_thread_child __bss setup_hpet disable_plane _idt_gate fgetc pdpte syscall_geral alloc_spin_lock hda_set_output_node sata_read_sector HDA_MEM free_frame idtr irq22 hda_inw keyboard_charset flush_tlb isr07 apic_timer irq7 speed task_switch set_ioapic_redir_table refresh_rate alloc_frame pit_set_frequencia fputc screen_refresh cmd_rename cmd_exit ioapic_cofiguration timer1 period pci_size call_function timer_wait setmsr lvt4 page_enable isr18 i2hex lvt_function ahci_initialize enable_NMI cmd_cd ap_startup pci_scan_bcc_scc setup_smp setup_hda irq0 fpu_save isr00 ata_initialize std_open_file std_putc rewind syscall_install syscall_writesector initialize_gui gdt_flush context_r13 isr06 lvt3 isr10 dv_num dsdt pipe_read mouse_y pci_scan_vendor syscall_tmpnam context_r10 cmd_echo syscall_alloc_pages lapicbase device_pde context_rip apic_timer_masked disable_NMI context_pid isr17 context_rbx enableapic hba_mem_space context_r14 irq21 ata_identify_device isr19 ret disable_pipe isr09 idt_flush isr30 strlen __code hda_outw filename_cmp clock ATA_BAR2 ATA_BAR5 read_super_block SLP_TYPb id_mouse_strings irq15 user_free timer3 acpi_virtual_addr cpuid_string gmbus_stoptransaction enable_dpll CORB_MEMORY g_mm_mp_index tss_install isr25 sata_idtfy ascii_maiusculas thread_setup context_rdi play_speaker setup_cursor KEYBOARD_BAT_TEST hda_max_volume HDBARU pci_write_config_dword ata_wait_no_drq cursor18x18 hda_send_verb gmbus_wait irq4 irq3 context_es input_node ioapic_masked  .symtab .strtab .shstrtab .text .data .got .got.plt .data.rel.local .bss .eh_frame .comment                                                                                     @             �                            !              �A      �      P                            '              �B      �     �                             ,             ��B     ��                                  5             ��B     ��     8                              E              C     �      4                             J              @E            0                             T      0                @     *                                                   0@     �G      
   
                	                       �     �                                                   ��     ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �b�  �����������                                                        ��   �� ��   ��  @�      ��1���f�X�  fg �f��"�ꐀ ��������������f� �؎������1�%�  ���  ������� ���� ������ ��1��� ���  �� ���$  �  � ���   � ���    0� ��%����� ���
   �����90  �����=�   t� ��� "��=0�  "߹�  �2   �    0 �   �"�� �  �p�   �������������H1��؎������H�% �  ��  �2�����0��  �2�  0H�%(�  �   ���H1��%8�  �    �H   "� �f���H��"��� �f���"�������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                Seja bem-vindo ao Sirius OS

	By: Nelson Cole
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ELF          >       �   @       h�         @ 8  @                   �      �                                      �      �   �        @                   P      ` �    ` �    0       0             Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��  ���_ cole _          �      �            � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           I��H�D �   L�H��C �   H�H�   �   L�H�  �   L�#H�  �   L�+�   �����H��H��H��H��L�������UH��AWSH��@��H�����I�      L�H�}�H�u�H�U�H�M�L�E�L�M�H���������H�H�U�H�H��     H�E�H�H�E�H�`     H�H�`     H�H� H��H��     H�H��     H�H��H�P     H�H�`     H�H�@H��H�H     H�H�E�H�h     H�H�E�H�@     H�H�E�H��     H�H��     H�H��H�X     H�I�߸    H��_������H���H�p     H�    H���������H�H� H��H�x     H�H���������H�H� H��H���������H�H� H�։�I��H���������H��ЉE�E��I��H�ú������H��АH��@[A_]���UH��AWSH����H�����I�%     L�H��j j�h  A�/ A��  �X  �   �d   H���������H�<I��H���������H���H�� H�E�H�E�H��I��H�T�������H���H���������H�H� �   H���r��   I��H���������H���H�E�H�E�H��������H�4H��I��H��r������H���H���������H�H� �   H�}�    �   I���rH�E�H��I��H�A������H�������UH��H��0��H�����I��     L�H�}�H�u��U܉M�L�E�H���������H�H� H�E��E�H9E�}?H�E��@��H9E�}0H�E�H�E��E�H�E�H��H�E�H�H��    H�E�HE؉������UH��SH��@��H�����I�`     Lۉ}ԉuЉỦM�L�E�L�M�f�E�  H�E�H�@H�E�H�E��@�E�}�u�E�    �E�    �   f�E� H�E��@�EȉE��H�H� H�E�H�� f�E�H�E�� ���E��J�E�f#E�f��t5�UЋE��Hc��UԋE��H�H�}��M�U�I��H��H���������H���f�e�m��}� y��E�H�E��@9E��b�����H��@[]���UH��AWSH��0��H�����I�I     Lۉ}܉u؉UԉM�D�E�L�M��E�    �X�E�    �CH�E�L��   �M�H�E��P�u؋E��Hc��}܋E��H�H��I��H���������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I��     Lۉ}܉u؉UԉM�D�E�L�M��E�    �p�E�    �[H�E�H��   �E��E�i��E��A��H�E��P�M؋E��Hc��M܋E��H�I��D��H��I��H���������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I��     Lۉ}܉u؉UԉM�D�E�L�M��}� �[  �}� �Q  �E�    �>H�E�L��   �M�H�E��P�E�Hc��}܋E��H�H��I��H���������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E����Hc��}܋E��H�H��I��H���������H��ЃE��E�;E�|��E�    �AH�E�H��   �M�H�E��P�u؋E��Hc��E�H�I��H��I��H���������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E��Hc��}܋E����H�H��I��H���������H��ЃE��E�;E�|���H��0[A_]���UH��AWSH��@��H�����I�)     Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}��  �E�    ��   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��   �E�f#E�f��tDH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H���������H����BH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H���������H���f�e�m��}� �[����E�H�E��@9E��	�����H��@[A_]���UH��SH��8��H�����I��     L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H���������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I�     Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}���   �E�    �   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��W�E�f#E�f��tBH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H���������H���f�e�m��}� y��E�H�E��@9E��T�����H��@[A_]���UH��SH��8��H�����I��     L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H���������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I�(     L�H�}ȉuĉU��M�D�E�D�M�H���������H�H� H�E�H�E�H   � �? �    H��I��H�p������H����E�    �U�H�E��P4�UH�E��P8�UH�E��P<H�E��@H   H�E��@L   H�E��P<H�E��PP�UH�E��PTH���������H�H��H�E�H�PXH�E��@D    H�E��PDH�E��P@�U�H�E��P�U�H�E��P�U�H�E��P �U�H�E��P�U H�E��P`�} u�E�   H�E��@�P�H�E��P(H�E��P�E�)ЍP�H�E��P$H�E��@0   �E����H�E��P,H�E��@��H�E��@��H�E�I���Ѻ    �    I��H�j�������H���H�E��@4��H�E��@����H�E�I��A�ȹ   �   �   H���������H��Ѓ}� u:H�E��@����H�E�I��A���� �   �   �   H���������H����8H�E��@����H�E�I��A���� �   �   �   H���������H��Ѓ}� t}H�E��@����H�U��E�I��A���� ����   �   H���������H���H�E��@4��H�E��@���ƋE��H�U�I��A�ȹ   ��ƿ   H���������H���H�E��@8A��H�E��@$��H�E��@(��H�E��@,��H�E��@0��H�E�I��H���������H���H�E�H��I��H�su������H������E�H�E�H�pHH�E��@��E܉������)Љ�H�E�H���u�I��A���� ������   ��H��H��������H���H��H�E��@����H�E�I��A�    �   �   �   H��������H���H�E�H�PHH�E��@��H���u�I��A���� ������   �ƿX   H���������H���H��H�E�H�PHH�E��@��(H���u�I��A���� ������   �ƿ-   H���������H���H��H�E�H�e�[A_]���UH��AWSH��0��H�����I��     L�H�}�H�u�H�E��P0H�E��@Ѓ�P�E�H�E��P,H�E��@Ѓ��E��E�P   �E�   �E�    �E���� H�E�H��I��H�su������H��ЉE�H�E�L�@H�M؋U܋E���������p��E�<�E��������ƋE���)ƋE��H�E�H���u�M��A�ȉщ�H��H�2�������H���H���H�e�[A_]���UH��H����H�����I��     L�H�}��   H�E�H���r�����UH��H����H�����I�g     L�H�}������UH��H����H�����I�<     L�H�}�H�U��BD    H�U��JDH�U��J@H�U��R8A��H�U��R$��H�U��R(A��H�U��R,��H�U��R0��H�U�I��D��I���������J��А����UH��SH��(��L�����I��     Mډ�f�E�H���������I�H� H�E�H���������I�H��H�E�H�PXH�E�@(�P�H�E�@H���к    ��E�H�E�@$�P�H�E�@L���к    ��E�H�E�P<H�E�PPH�E�PD�E�9�rH�E��@D    H�E�@@�PH�E�P@H�E�P@�E�9�r9H�E��@D    H�E�PDH�E�P@H�E�H��H���������I����E��  f�}���   H�E�@D����   H�E�@D�P�H�E�PDH�E�H�xHH�E�pTH�E�@PH�U�J,H�U�RLA��H�U�R@A��ʃ���H�U�J0H�U�RHA��H�U�RDA��ʃ�A��H���u�I��A������D�޿    H���������I���H����   f�}�	uH�E�@D�PH�E�PD��   f�}�
u!H�E��@D    H�E�@@�PH�E�P@�   f�}���   H�E�H�xHH�E�pTH�E�PPH�E�H,H�E�@LA��H�E�@@A��ȃ���H�E�H0H�E�@HA��H�E�@DA��ȃ�A���E�H���u�I��A���щ�D�މ�H���������I���H��H�E�@D�PH�E�PD�E�H�]�����UH��H����H�����I��
     L؉}�H���������H�H� H�E��U�H�E��P<�����UH��SH��(��H�����I��
     L�H�}�H�}� t=H�E�H�E��&H�E�H�PH�U�� f�����H�E�������H���H�E�� ��u���H��([]���UH��AWSH��P��H�����I�(
     L�H�}��u��U��M�L�E�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H��������H�<I�߸    H�Ϟ������H��Ҹ�����6  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H��������H�<I�߸    H�Ϟ������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�4�������H�<I�߸    H�Ϟ������H��Ҹ   ��   �E�    �   �E�    �   �}� tNH�E�H��   H�E��P�M��E���E��Hc��M��E���E��H��M�I��H��I��H���������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H���������H��ЃE��}� �U����E��}� �;����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��P��H�����I�F     L�H�}��u��U��M�D�E�L�M�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H��������H�<I�߸    H�Ϟ������H��Ҹ�����3  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H��������H�<I�߸    H�Ϟ������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�4�������H�<I�߸    H�Ϟ������H��Ҹ   ��   �E�    �   �E�    �   �}� tKH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H���������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H���������H��ЃE��}� �X����E��}� �>����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��0��H�����I�c     Lۉ}܉u؉U�H�M��E�    �   �E�    �t�U�������E��H���������H�Hڋ��E�}� tBH�E�H��   H�EȋP�MԋE��Hc��M؋E��H��M�I��H��I��H���������H��ЃE��}�~��E��}��o�����H��0[A_]���UH��AWSH��@��H�����I��     Lۉ}̉uȉUĉM�L�E��E���� �E�``` �E���� �EĉE��ẺE܋E��E؋EȉEԋE؍P��E��xH�M��E�I��A�    �   ��I��H��������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H��������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H��������H��ЋEԍP��E܍pH�M��E�I��A�    �Ѻ   ��I��H��������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H��������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H��������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H��������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H��������H��ЋEԍP��E܍p�M��E�ȃ�H�M�I��A�    �Ѻ   ��I��H��������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H��������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H��������H��ЋE؍P��M܋E�ȍp��E���H�M�I��A�    �   ��I��H��������H��АH��@[A_]���UH��AWSH��0��H�����I�U      Lۉ}܉u؉UԉM�D�E�D�M�H�} u
�    ��  �H   I��H���������H���H�E�H�}� u
�    ��  H�E�H   �    H��I��H�p������H���H�UH�E�H�P@H�E�U�PH�E�P0�E��H�E�PH�E�P,�E��H�E�PH�E��    H�E�P(�E�9�wH�E�P(H�E�P�
�U�H�E�PH�E�P$�E�9�wH�E�P$H�E�P�
�U�H�E�P�U�H�E�P�U�H�E�P H�E��@0    H�E�@0��I��H���������H���H��H�E�H�P8H�E�H�@8H��t.H�E�@0H�U�H�R8H�щ¾    H��I��H�p������H���H�E�@ ��H�E�@��H�E�@��H�E�@��H�E�@L�MA����I��H���������H���H�E�@��H�E�@��H�E�@��H�E�@L�MA�������I��H��������H���H�E�H��0[A_]���UH��AWSH�� ��H�����I��      L�H�}�H�E�H�@@H�E�H�E؋@ A��H�E؋@��H�E؋@��H�E؋@��H�E؋@��H�E�I��I��H���������H���H�E�H��H�>������H��АH�� [A_]���UH��AWSH�� ��H�����I�r�      L�H�}�H�}� u
������z  I�߸    H�-������H��҉E�}���   I�߸    H�-������H��҉E�}�[��   I�߸    H�-������H��҉E�}�Ct�}�Dt'�GH�E؋P,H�E؋@49�s1H�E؋@,�PH�E؉P,�H�E؋@,��tH�E؋@,�P�H�E؉P,����H�E�H��H�>������H��и    �  H�E�H�P8H�E؋@,��H�H�E��}� �C  H�E؋P,H�E؋@09��-  H�E��@    �}���   H�E؋@4��tkH�E؋@,��t`H�m�H�E؋P4H�E؋@,)�H�E�H�HH�E�H��H��I��H�?}������H���H�E؋@,�P�H�E؉P,H�E؋@4�P�H�E؉P4�   H�E��@   �~H�E؋P,H�E؋@49�t4H�E؋P4H�E؋@,)�H�E�H�HH�E�H��H��I��H�?}������H��ЋE��H�E��H�E؋@,�PH�E؉P,H�E؋@4�PH�E؉P4H�E��@   H�E�H��H�>������H���H�E؋@����u*H�E�H��H�>������H���H�E؋@����H�E؉P�    H�� [A_]���UH��AWSH��@��H�����I���      L�H�}�H�E�H�@@H�E�H�E�H�@8H�E��E�    f�E�  H�E��@��uH�E��@    �  �E�    �  �E�    �E�    ��   �}� ueH�E��P4�E�9�vH�E�H�PH�U�� f�f�E��f�E�  f�}�
uf�E�  �E�   H�E��P,�E�9�u�U�H�E��P$�U�H�E��P(�E�f�}� teH�E�H�xHH�E��p H�E��PH�E��H�E��A��H�E��H�E��A���E�H���u�I��A����D��D�։�I��H���������H���H���E�H�E��P�E�9������E�H�E��P�E�9������H�E�H�xHH�E��p H�E��@H�U��JH�U��R(�A��H�U��JH�U��R$�A��H���u�I��A����D��D�ֿ_   I��H���������H���H��H�e�[A_]���UH��AWSH��@��H�����I���      L�H�}�H�E��@ �E�H�E��@�E�H�E��@�E�H�E��@�E�H���������H�H� � �E�H���������H�H� �@�E�H���������H�H� �@�E̋EЃ����X  �E�;E�~Q�E���9E�~F�U�E��9E�}9�E��P�E��9E�})�E�+E��E�+E�։�I��H��������H�����   �E�;E���   �E�;E���   �U�E��9E���   �U��E��9E���   H���������H�H� � ��H�E��@ )ЉE�H���������H�H� �@��H�E��@)ЉE��aH���������H�H� � +EȉE�H���������H�H� �@+EĉE�}� y�E�    �}� y�E�    �U�H�E��P �U�H�E��PH���������H�H� �@����u�I�߸    H��������H��ҐH��@[A_]���UH��AWSH��@��H�����I���      L�H�}�H�u�H�UȉM�D�E�D�M��P  I��H���������H���H�E�H�E�P  �    H��I��H�p������H���H�E�H��I��H�su������H��ЉE�}�~�E�   �U�H�E�H�H0H�E�H��H��I��H��o������H���H�E��    H�E��U�P�U�H�E��P�E�����H�E��P�U�H�E��P�UH�E��PH�U�H�E�H�P(H�E�H�PHH�E��@����H�E��@����H�E�H��0H���u�I��A���� �    ��H��I��H�2�������H���H��H�E�H�U�H��H�e�[A_]���UH��AWSH��0��H�����I��      L�H�}�H�uЉU�H�E؋@$��H��H��H�H��H�PPH�E�H�H��H�E�H�E؋@$�HH�U؉J$H�U؉�H��H��H�H��H�H�PP�ẺH�E�H��I��H�su������H��ЉE�}�~�E�   �U�H�M�H�E�H��H��I��H��o������H��и    H��0[A_]���UH��AWSH��P��H�����I�%�      L�H�}��E�    �E�����H�E�H�@(H�E�H�E�H�PHH�E��@����H�E��@����H�E�H��0H���u�I��A���� �  � ��H��I��H�2�������H���H��H�E�H�PHH�E��@����H�E��@��H���u�I��A���� �  � ���H�N�������H�<I��H��������H���H��H�E؋P0H�E��@ЉE�H�E؋@,�E��E�d   �E�   �EĀ�� �E�    �H���������H�H� �@����u�H�E��@$���A  H�E��P$�E���A��H�}؋MċŰuЋE�I��A��D�щ�I��H���������H����E�    �  H���������H�H� � ��H�E؋@ )ЉE�H���������H�H� �@��H�E؋@)ЉE�H���������H�H� �@�E�E�Hc�H��H��H�H��H�PPH�E�H�H��H�E��E�;E���   �E��E��E�Ѓ�9E���   �UԋE��9E�}�E��E��E�E��9E�}gH�E�H�xH�MċE��E��E�ЍP�EԍpH�E�H���u�I��A�ȹ����H��I��H�2�������H���H���E��E�m��E����tZ�nH�E�H�xH�MċE��E��E�ЍP�EԍpH�E�H���u�I��A�ȹ    H��I��H�2�������H���H���E������E�H�E��P$�E�9��[����E�����A����}��t5H�M��E�Hc�H��H��H�H��H�H��P� ��I��H��������H����E�   �H���������H�H� �@����u�H�E�H�PHH�E��@����H�E��@����H�E�H��0H���u�I��A���� �    ��H��I��H�2�������H���H���E�H�e�[A_]���UH��AWSH����H�����I��      L�H�}�H�P       H�    H�X       H�    I�߸    H�[������H���H�`       �    H�}� t'H�E� ��H�`       �H�X       H�E�H��    H��[A_]���UH��AWH����H�����I�V�      L�H�`       �����   ����   ��t
��tA�   H�X       H�H����   H�X       H�H��I��H�������H����yH�X       H�H��tbH�S�������H�<I�׸    H�Ϟ������H����?H�X       H�H��t+H�X       H�H��I��H��#������H����������    H��A_]���UH��AWSH��@��H�����I�?�      Lۉ}��u�H���������H�H� H��t�}� x�}� y&�H���������H�H� �@����u������#  H�E�    H�E�    �E�    �E�    �E�    �E�    �   H��     �E�H�H�H��H�E�H�E�H��� �E�H�E�H��� �E�H�E�H��� �E�H�E�H��� �EċEԉE܋E�;E�~"�E�;E�~�UЋE��9E�}�ŰE��9E�|&�E��E�Hc�H���������H�H� H9��^������E�Hc�H���������H�H� H9�u&�H���������H�H� �@����u������  H�E� ���V  ����  ����  ���n  ��t����   �[  H��     �E�H�H�H��H��H�P       H�H�P       H�H�@(H�E�H�P       H��@��I��H��������H���H�P       H�H��I��H��������H��ЉE���  H��     �E�H�H�H��H��H�X       H�H�X       H�H�@@H�E�H�X       H��@��I��H��������H����E�    H�`       �   �H���������H�H� �@����u��]  H��     �E�H�H�H��H��H�X       H�H�X       H�H�@@H�E�H�X       H��@��I��H��������H����E�    H�`       �   �H���������H�H� �@����u���   H��     �E�H�H�H��H��H�X       H�H�X       H�H�@@H�E�H�X       H��@��I��H��������H����E�    H�`       �   �H���������H�H� �@����u��*�H���������H�H� �@����u��E�    ������I�}� t>��H�E�� ��u�H�E�� �PH�E��H�E�H��H�3������H���H�E��     �    H��@[A_]���UH��AWSH����H�����I���      L�H�}�H���������H�H� H��u*�   �    H��     H�<I��H�p������H���H���������H�H� H=�   ~�    �LH���������H�H� H�HH���������H�H�
H�U�H��     H�H��H���������H�H� H��[A_]���UH��AWSH�� ��H�����I���      L�H�}�H�E�    H�E؋@8A��H�E؋@$��H�E؋@(��H�E؋@,��H�E؋@0��H�E�I��I��H���������H����E�    �   H��     �E�H�H�H��H�E�H�E�� ��tWH�E�� ��uOH��     �E�H�H�H��H��H�X       H�H�X       H�H��I��H��������H��������E��E�Hc�H���������H�H� H9��\�����H�� [A_]���UH��AWSH�� ��H�����I���      Lۉ}�H�u�H�E�H��I��H�A������H��и    H��������H��҉E�E�H�� [A_]���UH��H����H�����I�!�      L؉}�H��     ���	v5H��     �D    H��     �    H��     �D    H��     ��JH��     �0�M�H��     ��H�0�L�H��     �T�JH��     �L�����UH��H����H�����I�]�      L�H��     �T��u
�    �   H��     �T��	vH��     �D    H��     �LH��     ��HT��U�H��     �T�JH��     �L0H��     ��H��D�    �E�����UH����H�����I���      L�H��     �D    H��     �    H��     �D    �]���UH��AWSH��0��H�����I�>�      L�H�}�H�u�H�E�H�E�H�Eȋ@��-�   �E�H�Eȋ@���2�E��E�,  �E�d   �EԍH��E؍P��E܍p�E���H�}�I��A�  ��I��H���������H��ЋEԍH��E؍P��E܍p�E���H�}�I��A�������I��H��������H���H�}ȋMԋU؋u܋E�I��A�������I��H��������H���H�E�H�HH�E܍P�E���
H���u�I��A�    �������H�Y�������H�<I��H��������H���H���E��E��m��m�J�EԍH��E؍P��E܍p�E���H�}�I��A�������I��H���������H��ЋEԍH��E؍P��E܍p�E���H�}�I��A�������I��H��������H���H�}ȋMԋU؋u܋E�I��A�������I��H��������H����E�    I�߸    H�-������H���f�E�f�}�
��   f�}� tl�}� ~ff�}�u_�m�f�E�  H�E�H�xH�E܍P�E��H�E����4�E�H���u�I��A������    ��I��H���������H���H��H�m��of�}� �\���H�E�H�xH�E܍P�E��H�E����4�E�H���u�I��A������    ��I��H���������H���H���E�H�E�H�PH�U��U҈������H�E��  ��H�Eȋ ��u�H�Eȋ �PH�EȉH�E�H��I��H�3������H���H�E��     �    H�e�[A_]���UH��AWSH��0��H�����I���      L�H�}��E���� �E�``` �E���� H�Eȋ@0��(�E�H�Eȋ@,��d�E��E�d   �E�2   �E؍P��E��xH�MȋE�I��A�    �   ��I��H��������H��ЋE؍P��E܍p�E���H�}ȋM�I��A�ȹ   ��I��H��������H��ЋE؍P��E܍p�E���H�}ȋM�I��A�ȹ   ��I��H��������H��ЋEԍP��E܍pH�MȋE�I��A�    �Ѻ   ��I��H��������H��ЋEԍP��E܍p�E���H�}ȋM�I��A�ȉѺ   ��I��H��������H��ЋEԍP��E܍p�E���H�}ȋM�I��A�ȉѺ   ��I��H��������H��ЋEԍP��E܍p�M��E�ȃ�H�}ȋM�I��A�ȉѺ   ��I��H��������H��ЋEԍP��E܍p�M��E�ȃ�H�}ȋM�I��A�ȉѺ   ��I��H��������H��ЋEԍP��E܍p�M��E�ȃ�H�M�I��A�    �Ѻ   ��I��H��������H��ЋE؍P��M܋E�ȍp��E���H�}ȋM�I��A�ȹ   ��I��H��������H��ЋE؍P��M܋E�ȍp��E���H�}ȋM�I��A�ȹ   ��I��H��������H��ЋE؍P��M܋E�ȍp��E���H�M�I��A�    �   ��I��H��������H��АH��0[A_]���UH��AWSH��0��H�����I���      Lۉ}܉u؉UԉM�D�E�D�M�H�} u
�    ��  �H   I��H���������H���H�E�H�}� u
�    ��  H�E�H   �    H��I��H�p������H���H�UH�E�H�P@H�E�U�PH�E�P0�E��H�E�PH�E�P,�E��H�E�PH�E��    H�E�P(�E�9�wH�E�P(H�E�P�
�U�H�E�PH�E�P$�E�9�wH�E�P$H�E�P�
�U�H�E�P�U�H�E�P�U�H�E�P H�E��@0    H�E�@0��I��H���������H���H��H�E�H�P8H�E�H�@8H��t.H�E�@0H�U�H�R8H�щ¾    H��I��H�p������H���H�E�@ ��H�E�@��H�E�@��H�E�@��H�E�@L�MA����I��H���������H���H�E�@��H�E�@��H�E�@��H�E�@L�MA�������I��H��������H���H�E�H��0[A_]���UH��AWSH��0��H�����I�X�      L�H�}�H�}� u
������,  I�߸    H�-������H��҉E�}���   I�߸    H�-������H��҉E�}�[uqI�߸    H�-������H��҉E�}�At�}�Bt �2H�Eȋ@,��t&H�Eȋ@,�P�H�EȉP,�H�Eȋ@,�PH�EȉP,��H�E�H��H�
%������H��и    �pH�E�H��I��H�W�������H���H�E�H�EȋP(H�E�� 9�s=H�E�� ��H�EȉP(H�Eȋ@(��:vH�E��@(    H�E�H��H�
%������H��и    H��0[A_]���UH��AWSH��@��H�����I���      L�H�}�H�E�H�@@H�E�H�E�H�@8H�E�H�E�@   H��H�t�������H�<I��H�SQ������H��ЉE��E�    H�E��@���E���H�EЋ ��u�H�EЋ �PH�EЉ�E�    �!  H�E��@�E�H�E��@ �E�H�E��P,�E�9�u�E�i� �E�����H�E��@��A��H�E��@�U���Ѓ���H�E��@����H�UЋE�I��A���   D��I��H���������H��ЋE�;E���  H�E�H��H��'������H���H�E�H�xH�u؋U�H�E��@�M���ȃ�A��H�E��H�E�ȃ�A��H�E�H���u�I��A����D��D��H��I��H��������H���H��H�E��@��E�ЉE�H�E�H�xH�u؋E�H�U��R�M���ʃ�A��H�U��J�U�ʃ�A��H���u�I��A����D��D��H�p       H�<I��H��������H���H��H�E��@���E�ЉE�H�E�H�xH�u؋E�H�U��R�M���ʃ�A��H�U��J�U�ʃ�A��H���u�I��A����D��D��H��       H�<I��H��������H���H���E�    H�m考E��E�;E������H�E��     �H�e�[A_]���UH��AWSH��@��H�����I���      L�H�}�H�E��@b���� ����  H�w�������H�H�|�������H�4H��       H�<I�߸    H��������H���H�E��@o��H��x�H*��H��H���H	��H*��X��E�H�����������E��E�    H�E��@o=���?v�E�   H�����������E��)H�E��@o=�� v�E�   H�����������E��E��^E��E�H�E�fHn�H��������H�4H�p       H�<I�߸   H��������H���H�p       H�<I��H�su������H��ЉE̋ẺE��H�p       �E�H�H�� �E��}�~�H�        �E�H�H�H��H�w       H�H�|�������H�4H��I�߸    H��������H����   H���������H�H�|�������H�4H��       H�<I�߸    H��������H���H���������H�H�|�������H�4H�p       H�<I�߸    H��������H��ѐH��@[A_]���UH��AWSH����H�����I�d�      Lۉ}�H�u�H�E�� ��H�E��@9�sH�E��P#H�E��@9�r"H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@��u)H���������H�H��E�H�։�H��*������H���H�E�H�PH�E��@#��H�H�E�H�PH�E�H�@�U�H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  H�E��@��u0H���������H�H� H��t�E�����I��H�E�������H��ЋE�H��[A_]���UH��H����H�����I��      L�H�}��E�    H�E�@��u]H�E�@'�PH�E�P'��H�E�P#H�E�@'9�r�H�E�H�PH�E�@'��H��H�H�E�H�PH�E�H�@� ���E��   H�E�@��tH�E�@��uiH�E�@#��u������ZH�E�P'H�E�@#9�r������AH�E�H�PH�E�@'��H�H�E�H�PH�E�H�@� ���E�H�E�@'�PH�E�P'�E�����UH��H����H�����I���      L�H���������H�H� H�E��E�    H�E��@��uWH�E��P#H�E��@'9�w�    �AH�E�H�PH�E��@'��H�H�E�H�PH�E�H�@� ���E�H�E��@'�PH�E��P'�E�����UH��H����H�����I�G�      L�H���������H�H� H�E��E�    H�E��@��uXH�E��@'�PH�E��P'��H�E��P#H�E��@'9�r�H�E�H�PH�E��@'��H��H�H�E�H�PH�E�H�@� ���E��E�����UH��AWH��(��H�����I���      L�H�}�H�u�H�U����u�    �(H�M�H�U�H��H��I��H�-F������H���H�E�H�E�H��(A_]���UH��AWSH�� ��H�����I�+�      L�H�}�H�}� u
������   H�}� tH�E؋@����tH�E��@"<t������zH�E؋@%�   ��u�    �cH�E؋@#H�U؋J�    ��E�H�E؋@��@��u�U�H�E؉�H��I��H�P������H���H�E�H��I��H�qM������H��ЉE�E�H�� [A_]���UH��AWSH����H�����I�D�      L�H�}�H�}� u������0H�E�H��H��.������H���H�E�H��I��H��N������H���H��[A_]���UH��AWSH�� ��H�����I���      Lۉ}�H�u�H�}� u
�������  H�EЋ@��u
�    �  H�EЋ@��tH�EЋ@��tH�EЋ@��u!H�UЋE�H�։�H��*������H����y  H�EЋ@����unH�EЋP#H�EЋ�+  9�wYH�EЋ�+  ��tKH�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��E�U�H�EЉ�H��I��H��O������H����H�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U܈H�E�� ��H�EЋ@��9�r3H�EЋ@����H�EЉPH�E�f�   H�E�H��H��.������H���H�EЋ@#�PH�EЉP#H�EЋP#H�EЋ�+  9�vH�EЋ�+  �PH�EЉ�+  H�EЋ@���H�EЉP�    H�� [A_]���UH��AWH��(��H�����I���      L�H�}�H�}� u
������  H�E؋@��u
�    �v  H�E؋@��tH�E؋@��tH�E؋@��u"H�E�H��H��+������H��ЉE�E��0  H�E؋P#H�E؋�+  9�r
������  H�E؋@����ulH�E؋P#H�E؋�+  9�wWH�E؋�+  ��tIH�E؋@����H�E؉PH�E؋@#H�U؋r�    ���E�U�H�E؉�H��I��H��O������H���H�E؋@#H�U؋J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@� ���E�H�E�� ��H�E؋@��9�rH�E؋@����H�E؉PH�E�f�   H�E؋@#�PH�E؉P#�E�H��(A_]���UH��SH��H��H�����I���      L�H�}ȉuĉU�H�M�H�}� u�    �y�E�    H�E�H�E��E�    �FH�E�H��H�;2������H��ЉE؃}��u�E�    �u��4H�E�H�PH�U��U؈�E��E��E��E��E�9�w��E�    �u�H��H[]���UH��SH��H��H�����I�(�      L�H�}ȉuĉU�H�M�H�}� u�    �l�E�    H�E�H�E��E�    �9H�E�H�PH�U�� ���E�H�U��E�H�։�H�0������H��ЃE��E��E��E��E�9�w��E�    �u�H��H[]���UH��H����H�����I�u�      L�H�}�H�u��U�}�tZ�}�|�}� t�}�t�nH�E���H�E��P#H�E���H�E��P'�RH�E��@#H�U��H�E��P#H�E��@'H�U��H�E��P'�(H�E���+  H�U�)Љ�H�E��P#H�E��P#H�E��P'�H�E��@#H�U��J�    ��Љ�H�E�f��    ����UH��H����H�����I���      L�H�}�H�}� u�    �	H�E��@#������UH��H����H�����I�V�      L�H�}�H�}� t7H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@����H�E��P������UH��H��(��H�����I���      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H��(��H�����I���      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H����H�����I�C�      L�H�}��E�_   �(�E�Hc�H�E�H�� < u�E�Hc�H�E�H��  �m��}� y����    ����UH��H����H�����I���      L�H�}�H�E�H�E�H�E�H�E��H�E�� </uH�E�H��H�E�H�E�H�E�� ��u�H�E�����UH��H��0  ��H�����I�p�      L�H������H������H������H�E�H������H�E�H������H�E��E�    �?H�E�� ��u�E�Hc�H�E�H��  �H�E�H�PH�U��U�Hc�H�U�H�� ��E��}�_~��E�    �-H�E�H�PH�U��H�E�H�PH�U�� 8�t�   ��E��}�_~͸    ����UH��SH�� ��H�����I���      L�H�}�H�u�H�E؋PH�E؋@ЉE�E�H�U����H�     H�H�¾   H�7������H��ЉE�}� t
�������   �E�    ��   �E�%�  ��H�     ��H؋���uf�E�%�  ��H�     ��H��������E�H�U����H�     H�H�¾   H�\7������H��ЉE�}� t������r�E��m�E�%�  =�  uE�E��E�H�U����H�     H�H�¾   H�7������H��ЉE�}� t�������E�H�E؋@$9E����������H�� []���UH��H����H�����I��      L؉}��u�H�U�H�M�    ����UH��AWSH��0��H�����I���      Lۉ}�H�u�H�U�H�EȋPH�Eȋ@ЉE�H�Eȋ@ �E܉E�ЉE�   �    H�     H�<I��H�p������H����E�    �B�U�E�Љ�H�EЋ ��H�     H��   H�\7������H��ЉE��}� u�E�H�EȋP �E�9�w���H��0[A_]���UH��H����H�����I���      L�H�}�H�u�H�U��R��H�U����H�U�H��H��   I�7������J� ������UH��AWSH��`��H�����I��      L�H�}�H�u�H�U�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�E�H�E�H�E�H��I��H��m������H��ЉE�H�E��@,�E��9  H�E�H�E��H�E�� </uH�E��  H�E��H�E�H�E�� ��u׋U�H�E��@ H�M��	��H�M���H�7������H��ЉE؃}� t#H�E�H��I��H� �������H��и    ��   �E�    �f�E���Hc�H�E�H�H�E�H�E��@a��t5H�E��@b����@��t#H�E�H�U�H��H��H��8������H��ЉE���E������}� t�E��}�?~����}� u+�}�?%H�EЋ@k�E�H�E��@ �E؉E�ЉE�m��	�E�    �
�}� �����H�E�H��I��H� �������H��ЋE�H��`[A_]���UH��AWSH��P��H�����I�j�      L�H�}�H�u�H�U��M�L�E�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�Eغ    �    H��I��H�p������H��ЋU�H�E��@ H�M��	��H�M؉�H�7������H��ЉE�}� t#H�E�H��I��H� �������H��и������   �E�    �T�E���Hc�H�E�H�H�E�H�E��@a��t#H�E�H�U�H��H��H��8������H��ЉE���E������}� t�E��}�?~����}� u:�}�?4�E���Hc�H�E�H�H�EȺ�   H��H��I��H��o������H�����E�����H�E�H��I��H� �������H��ЋE�H��P[A_]���UH��AWSH��P��H�����I���      L�H�}�H�u�H�U�H�E���C  ��u
������	  H�E���C  ��@v/H���������H�<I�߸    H�Ϟ������H��Ҹ������  H�E��PH�E��@ЉE�H�E���?  H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�Eغ    �    H��I��H�p������H��ЋU�H�E��@ H�M��	��H�M؉�H�7������H��ЉEԃ}� t!H�E�H��I��H� �������H��ЋE��  H�E���C  ��H��H��H�E�H�H�E�H�EȺ`   �    H��I��H�p������H���H�E�H��+H��H�8������H���H��H�E�H��H��I��H��r������H����E�    �"H�UȋE�H����uH�UȋE�H�� �E��}�_~�H�E��@` H�E���+  H�EȉPo�U�H�E��@ H�M��	��H�M؉�H�\7������H��ЉE�H�E�H��I��H� �������H��ЋE�H��P[A_]���UH��AWSH��`��H�����I�C�      L�H�}�H�u�H�U��S  I��H���������H���H�E�H�EкS  �    H��I��H�p������H���H�E��PH�E��@ ��H�EЉP�    I��H���������H���H�U�H�BH�E��PoH�EЉ�+  H�E��PH�EЉ�/  H�E��P H�EЉ�3  H�E��H�EЉ�G  �    I��H���������H���H�U�H��K  H�E�H��K  �    �    H��I��H�p������H���H�E��@k�E�    I��H���������H���H�E��E������E�    �E�    ��  �   I��H���������H���H�U�H��K  �M�Hc�H��H�H�H�E�H��K  �U�Hc�H��H�H� H�E�H�E��   �    H��I��H�p������H����E�    �<  H�E��@ �E��H�E��@�H�E��P�E�H�H�4�    H�E�H�ʉH�EЋ�;  �PH�EЉ�;  �E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E�;E�ts�E�H�U����H�U�H��H�¾   H�7������H��ЉE��}� t:H�E�H��I��H� �������H���H�E�H��H��N������H��и    �   �E��E�H�E��@�����E�    ��U�E�H��    H�E�HЋ �E�}��u	�E�������E��}��  ������}��t�E��}��  � �����H�E�H��I��H� �������H���H�E�H��`[A_]���UH��AWSH��p  ��H�����I���      L�H������H�������   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H������H�E�H��H��I��H�bk������H���H�U�H�E�H��H��I��H�n������H��п�   I��H���������H���H��     H�H��     H���   �    H��I��H�p������H��п   I��H���������H���H�E�H�EȺ   �    H��I��H�p������H���H�E�H�E�H�E��   �    H��I��H�p������H����E�    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ ���    Hǅ���    Hǅ���    Hǅ���    Hǅ ���    Hǅ(���    Hǅ0���    Hǅ8���    Hǅ@���    HǅH���    HǅP���    HǅX���    Hǅ`���    Hǅh���    Hǅp���    Hǅx���    H�E�    H�E�    H������H������H��H��I��H��r������H���������<wt������<au�E�   H�E��@   H�E��     H�U�H�E�H��H��H�<������H��ЉE�}� t_H��     H�H��I��H� �������H���H�E�H��I��H� �������H���H�E�H��I��H� �������H��и    �  H�E�H�U�H�M�H�E�H��H��H�r<������H��ЉE��}� u_H��     H�H��I��H� �������H���H�E�H��I��H� �������H���H�E�H��I��H� �������H��и    �  H�EȋU��P,H��     H�H�M�H�U�H�u�I�ȹ    H��H��>������H��ЉE�}����   �}� tqH��     H�H������H�U�H�u�A�    H��H�BU������H���H��     H�H������H�U�H�u�I�ȹ    H��H��>������H��ЉE�}� ��   H��     H�H��I��H� �������H���H�E�H��I��H� �������H���H�E�H��I��H� �������H��и    ��  �}� t_H�E�H��I��H� �������H���H��     H�H��I��H� �������H���H�E�H��I��H� �������H��и    �r  H��     H�H�U�H�M�H��H��H��B������H���H�E�H�}� ��   H��     H�H��H�E�H��+�`   H��H��I��H��o������H���H�E�H��+H��H��7������H���������<wt������<+t������<au
H�E��@"�H�E��@"H�E��@   H�EȋP,H�E���?  H��     H��PsH�E���C  ������<auH��     H��PoH�E��P#H�E�H��I��H� �������H���H��     H�H��I��H� �������H���H�E�H��I��H� �������H���H�E�H��p  [A_]���UH��AWSH��@��H�����I���      L�H�}��   I��H���������H���H�E�H�E�   �    H��I��H�p������H���H�E�H�E�H�E�   �    H��I��H�p������H���H�E��@   H�E��     H�U�H�E�H��H��H�<������H��ЉE܃}� t H�E�H��I��H� �������H��и�����AH�U�H�M�H�E�H��H��H�Q@������H��ЉE�H�E�H��I��H� �������H��ЋE�H��@[A_]���UH��AWSH�� ��H�����I�F�      L�H�}�H�E�H�@H��I��H� �������H����E�    �TH�E�H��K  �U�Hc�H��H�H� H��t?H�E�H��K  �U�Hc�H��H�H� H��I��H� �������H��ЃE��}��  ~���H�E�H��K  H��I��H� �������H���H�E�H��I��H� �������H���H�E�    �    H�� [A_]���UH��H�� ��L�����I�I�      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H�7������I� ������UH��H�� ��L�����I�u�      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H�\7������I� ������UH��AWSH��   ��H�����I���      L�H��x���H��p�����l����   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H��x���H�E�H��H��I��H�bk������H���H�U�H�E�H��H��I��H�n������H��п   I��H���������H���H�E�H�EȺ   �    H��I��H�p������H���H�E�H�E�H�E��   �    H��I��H�p������H���H�E��@   H�E��     H�U�H�E�H��H��H�<������H��ЉE��}� t_H��     H�H��I��H� �������H���H�E�H��I��H� �������H���H�E�H��I��H� �������H��и�����-  H�E�H�U�H�M�H�E�H��H��H�r<������H��ЉE��}� u_H��     H�H��I��H� �������H���H�E�H��I��H� �������H���H�E�H��I��H� �������H��и�����  H�EȋU��P,H�EȋPH�Eȋ@ЉE�H�EȋP,H�Eȋ@ �ЋE�ЉE��    I��H���������H���H�E�H�E��    �    H��I��H�p������H��ЋU�H�Eȋ@ H�M��	��H�M���H�7������H��ЉE��E�    �E�    �   �E���Hc�H�E�H�H�E��E�;�l���}~H�E��@a��ta�E���Hc�H��p���H�H�E���   H��H��I��H��o������H��ЋE���Hc�H��p���H�H��H��7������H��ЃE����E��}�?�e�����H�E�H��I��H� �������H���H�E�H��I��H� �������H���H�E�H��I��H� �������H��ЋE�H�Đ   [A_]���UH��AWSH��`��H�����I���      L�H�}�H�u�H�U�H�M�D�E�H�E�H�E�H�Eغ�   �    H��I��H�p������H���H�E�H��H�8������H���H��H�E�H��H��I��H��r������H����E�    �"H�U؋E�H����uH�U؋E�H�� �E��}�_~�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉEп    I��H���������H���H�E�H�EȺ    �    H��I��H�p������H��ЋU�H�E��@ H�M��	��H�Mȉ�H�7������H��ЉEă}� t!H�E�H��I��H� �������H��ЋE���  �E�    �$�E���Hc�H�E�H�H�E�H�E��@a��t�E��}�?~���H�E��@a���G  �}�?�=  �U�H�E؉PsH�E��@a��E���H�E؈PbH�U�H�E�H��H��H�h9������H���H�U؉BkH�E؋@k���uOH�E�H��H���������H�<I�߸    H�Ϟ������H���H�E�H��I��H� �������H��и   ��   �E���@��t$H�E؋@kH�U�H�M�H�Ή�H�+;������H���H�M�H�E຀   H��H��I��H��o������H��ЋU�H�E��@ H�M��	��H�Mȉ�H�\7������H��ЉEĐH�E�H��I��H� �������H��и    �JH�E�H��I��H� �������H���H�E�H��H���������H�<I�߸    H�Ϟ������H��Ҹ����H��`[A_]���UH��AWSH��P��H�����I�F�      Lۉ}�H�u�H�U��    I��H���������H���H�E��E�    �E��E��E������E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E��E܋E�;E���   �}� tV�E�H�U����H�U�H��H�¾   H�\7������H��ЉẼ}� t#H�E�H��I��H� �������H��и�����?  �E�H�U����H�U�H��H�¾   H�7������H��ЉẼ}� t#H�E�H��I��H� �������H��и������   �E��E�E��E��E�   H�E��@�����E�    ��U�E�EȋE�H��    H�E�HЋ �E�E�H��    H�E�H��     �}��uL�E�H�U����H�U�H��H�¾   H�\7������H��ЉE̐H�E�H��I��H� �������H��ЋE��6�E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��Y���H��P[A_]���UH��AWSH��   ��H�����I���      L�H��h����   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H��h���H�E�H��H��I��H�bk������H���H�U�H�E�H��H��I��H�n������H��п   I��H���������H���H�E�H�E��   �    H��I��H�p������H���H��p���H�E�H�E��   �    H��I��H�p������H���H�E��@   H�E��     H�U�H�E�H��H��H�<������H��ЉE�}� t<H�E�H��I��H� �������H���H�E�H��I��H� �������H��и    ��  H�E�H�U�H�M�H�E�H��H��H�r<������H��ЉE��}� u<H�E�H��I��H� �������H���H�E�H��I��H� �������H��и�����d  H�E��U��P,H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE��    I��H���������H���H�E�H�E��    �    H��I��H�p������H��ЋU�H�E��@ H�M��	��H�M���H�7������H��ЉE�}� tSH�E�H��I��H� �������H���H�E�H��I��H� �������H���H�E�H��I��H� �������H��ЋE��l  �E�    �   �E������E���Hc�H�E�H�H�E�H�E��@a��t!H�E�H�U�H��H��H��8������H��ЉE�}� u9H�E��@a �U�H�E��@ H�M��	��H�M���H�\7������H��ЉE�}� ��E��}�?�k����}� tPH�E�H��I��H� �������H���H�E�H��I��H� �������H���H�E�H��I��H� �������H��ЋE��uH�E��@kH�U�H�M�H�Ή�H��X������H��ЉE�H�E�H��I��H� �������H���H�E�H��I��H� �������H���H�E�H��I��H� �������H��ЋE�H�Đ   [A_]���UH��H����H�5����I���      Lމ}�E�E��}� u�E��   �E����rH�      H�H�      H�����UH��H����H�����I�;�      L�H�}��   H�E�H���r�����UH��AWH����H�����I� �      L�H�     H�H�U�H�     H�    H��       �    H�M�   �    H��I��H�p������H��ѐH��A_]���UH��AWSH��P��H�����I�x�      Lۉ}��u��}� u
�    ��  H�     H�H=�   v%H�8�������H�<I�߸    H�Ϟ������H��ҐH��       ���u�H��       ��PH��       ��E����E�E�%�  ��t�E��E�    �E�    �E�    �}� t�E��   �E�   �K  �}��  �=  H�     H�H�E�H�E�    �E�    �  H�E؋@����   H�E؋@9E���   H�E�H�H�E؋@��H�H�E�H�E؋@+E���H�E؉PH�E؋P�E��H�E؉PH�E�H�E�H�     H�H�E��E�    �mH�E؋@��tH�E��E��WH�E�H�E�H�E�H�E�H�E�H�@H�PH�E�H�PH�E��@   H�E�H�U�H�H�E��U��PH�E�H�U�H�P�E���!�}��   ~��H�E��E��}��   ������E�   ���}� ��   H�     H�H�E��E�    �~H�E؋@��tH�E��E��hH�E�H�E��E��H�X_������H���H�E�H�E�H�U�H��E��E���H�E��PH�E��U��P�E���+E���H�E��PH�E�H�@   ��}��   �u���H��       �    H�     H�H�PH�     H�H�E�H��P[A_]���UH��SH��(��H�����I�S�      L�H�}�H�}� ��  �H��       ���u�H��       ��PH��       �H�E�H�E�H�     H�H�E��E�    �M  H�E�H� H9E�tH�E��E��2  H�E�H�E�H�     H�H�P�H�     H�H�E؋@��uH�E�H��H��_������H����   H�E؋@��uH�E�H�@H�E�H�E�H�@H�P�H�E�H�PH�E�H�@H��tH�E؋@����   H�E�H�@H��uRH�E�H� H��H��_������H���H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    ��}��   �������H��       �    ��H��([]���UH��AWH��H��L�����I�Q�      M�H�}��u�H�E�    �E�    H�}� u�E��   ��H�y`������I� ���8  �H��       A� ��u�H��       A� �PH��       A� H�     I� H�E�H�E�H�E��E�    �   H�E�H� H9E�t
H�E��   H�E�H�E��E�   H�E��P�E��=   v@H�     I� �U�H�E�H��H�p�������I�< M�Ǹ    I�Ϟ������M�A����H�E�H� H�E�H�E��P�E��H�E��P�E��}��   �X���H��       A�     �}� u�E��   ��H�y`������I� ���H�E�H��HA_]���UH��H�� ��H�����I���      L�H�}�H�u��E�    H�E�H�E��   H�E�� ��H�E��@9�sH�E��P#H�E��@9�rH�E��@#    H�E�f�   H�E�H�PH�E��@#��H�H�E�H�PH�E�H�PH�U�H�U�H�R� �H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  �E��}��E����E�����UH��H�� ��H�����I���      L�H�}�H�u��E�    H�E�H�E�H�E��@'�PH�E��P'H�E��P'H�E��@9�rH�E��@'   �H�E��P#H�E��@'9�r�H�E��@'�P�H�E��P'�JH�E�H�PH�E��@'��H�H�E�H�PH�E�H�PH�E�H�HH�M���H�E��@'�PH�E��P'�E��}�~��E�����UH��AWSH��0��H�����I�ʖ      L�H�}�H���������H�H� H�E�H�E�H�E�H�E�H��I��H�su������H��ЉE�H�E�H��I��H�su������H��ЉE؋U܋E��=   ~
������   H�E�� </uH�E��E�H�HE�H�m�H�E�� </tH�E�H�E�H�PH�U�� /�H�E�H�U�H�E�H��H��I��H��r������H���H�E�H��I��H�su������H��Љ�HE�H�m�H�E�� </u	H�E��  �H�E�H�E��  �    H��0[A_]���UH��AWSH����H�����I�{�      L�H���������H�H� H��I��H�su������H��Ѓ�w
�    �   H���������H�H� H�E�H�E�H��I��H�su������H��Љ�HE��H�E�H�P�H�U��  H�E�� </u�H���������H�H� H��I��H�su������H��Ѓ�vH�E��  �    H��[A_]���UH��AWSH��0��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
�    ��  H�E�H��I��H�su������H��ЉE�E�H�H�P�H�E�H�� </u�E�H�H�P�H�E�H��  �}� 
�    �  �}���   H�E�H��� <:u%H�U�H�E�H��H��I��H��r������H����K  H���������H�<I��H���������H���H��H�E�H��H��I��H��r������H���H�E�H��I��H�su������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H��r������H����   H���������H�<I��H���������H���H��H�E�H��H��I��H��r������H���H�E�H��I��H�su������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H��r������H���H�E�H��0[A_]���UH��H����H�����I�O�      L�H�}�H�E�H�E�H�}� u�    �+�E�    �H�E�� </u�E�H�E�H�E�� ��u�E�����UH��AWSH��0��H�����I��      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
������   H�E�H��I��H�su������H��ЉE�E�H�HE�H�m��H�E�� </tH�m�H�E�� ��t�E�P��U�����H�E�H�U�H�E�H��H��I��H��r������H���H�E��  �    H��0[A_]���UH��H��8��H�����I���      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �CH�E�H�PH�U�� ���E�H�E�H�PH�U�� ���E�E�+E�E�}� u�}� t
�m��}� u��E�����UH��H��8��H�����I�f�      L�H�}�H�uЉŰẺE�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M����E��P��U���u�H�E�����UH��H�� ��H�����I��      L�H�}���U��E�E��E�H�E�H�E��H�E�H�PH�U��U��m��}� u�H�E�����UH��AWSH��0��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E��E�    H�E�H�PH�U�� ����I��H��~������H��ЉE�H�E�H�PH�U�� ����I��H��~������H��ЉEԋE�+EԉE܃}� u�}� t뗋E�H��0[A_]���UH��AWSH����H�����I�ώ      L�H�}�H�u�H�E�H��I��H�su������H��Љ�H�E�H�H�E�H��H��I��H��r������H���H�E�H��[A_]���UH��H�� ��H�����I�X�      L�H�}�u�H�E�H�E��H�E�� ��9E�uH�E��H�E�H�E�� ��u۸    ����UH��H�� ��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E��3H�E��H�E�� 8�u!H�E�� ��H�E�� ��Ѕ�u�    �'H�E�H�PH�U��H�E�H�PH�U�� 8�t����������UH��H��0��H�����I�]�      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E��  H�E�����UH��AWH��(��H�����I���      L�H�}؉uԋU��҉Uԃ}� uOH�U�H��I��H�su������H��҉�H�E�H���   H�E�� ��tH�E�� ��9E�u	H�E��   H�E�H�E؃�H��űE�i��E�H�E�H�E��H�E�H�E� ������H�E� ��!�%������u%H�E� 3E䍐����H�E� 3E���!�%������t�H�E�H�E��H�E�H�E�� ��tH�E�� ��9E�u�H�E�H��(A_]���UH��H��@��H�����I���      L�H�}�H�u�H�U�H�U�H�U������   H�U�H�������   H�E�    H�E�    H�E�    H�E�    �H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�t�H�E�H+E��'H�U����H�Uȉ�H��H�s������H���H+E�����UH��H����H�����I���      L�H�}�H�E�H�E��H�E�H�E�� ��u�H�E�H+E�����UH��AWSH��@��H�����I�2�      L�H�}�H�u��U�H�E�H�E�H�E�H�E��E�    �kH�E�H�PH�U�� ����I��H��~������H��ЉE�H�E�H�PH�U�� ����I��H��~������H��ЉEԋE�+EԉE܃}� u�}� t
�m��}� u��E�H��@[A_]���UH��H��(��H�����I�m�      L�H�}�H�u��U�H�E�H�E�H�E�H�E��}� u)������2H�E�H�PH�U��H�E�H�PH�U�� 8�u�m��}� u����E�����UH��H��8��H�����I��      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �!H�U�H�BH�E�H�E�H�HH�M����E��E�9E�w�H�E��  �E�����UH��AWH����H�����I�n�      L�H�}�H�u�H�M�H�U�H��H��I��H�=t������H��҉�HE�H�E�� ��tH�E���    H��A_]���UH��AWH��(��H�����I���      L�H�}؉u�H�U�H��I��H�su������H��҉E��U�H�E�H�H�E��E�    �H�E�� ��9E�uH�E��H�m��E��E�9E�wڸ    H��(A_]���UH��H��0��H�����I�k�      L�H�}�H�u�H�E�H� H�E�H�}� u�    �vH�E�H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u,�}� u
H�E�    �H�E�H���  H�E�H�U�H�H�E���}� u������UH��H��@��H�����I���      L�H�}�H�u�H�E�H�E�H�E�    H�E�    H�E�    H�E�    H�E�� ��u
�    ��   H�E�H��� ��u+�H�E�H�E��H�E�� 8�t�H�E�H+E��   H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�u�H�E�H+E�����UH��H��8��H�����I�{�      L�H�}�H�u�H�U�H�}� uH�E�H� H�E�H�}� u
�    ��   �H�E�H�PH�U�� ���E�H�E�H�E��
�E�;E�u��H�E�H�PH�U�� ���E��}� uۃ}� uH�E�H�     �    �   H�E�H��H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u4�}� u
H�E�    �H�E�H��H�E�H�E��  H�E�H�U�H�H�E���}� u������UH��H����H�����I�D�      L�H�}�H�u�H�u�H�M�H��       H�H��H�yz������H�������UH��AWSH�� ��H�����I��      L�H�}�H�u�H�E�H��I��H�su������H��ЉE��2�U�H�M�H�E�H��H��I��H��n������H��Ѕ�uH�E��H�E�H�E�� ��uø    H�� [A_]���UH��AWSH�� ��H�����I�R�      L�H�}�H�E�H��I��H�su������H��Ѓ��E�E��I��H���������H���H�E�H�}� u�    �$�U�H�M�H�E�H��H��I��H��o������H��АH�� [A_]���UH��H��8��H�����I���      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��U�H�E�H�H�E�H�E�H;E�v[H�E�H;E�sQH�E�H�E��E�HE��H�m�H�m�H�E��H�E��H�E�H;E�u��'H�U�H�BH�E�H�E�H�HH�M���H�E�H;E�u�H�E�����UH��AWH����H�����I��      L�H�}�H�u�H�M�H�U�H��H��I��H��q������H���H��A_]���UH��AWH����H�����I���      Lډ}�H���������H�<I�׸    H�Ϟ������H�������UH��H����H�����I�M�      L؉}��U���H���������H�Hc��������t�E� �E�����UH��H����H�����I���      L؉}��U���H���������H�Hc��������t�m� �E�����UH��AWSH��0��H�����I���      L�H�}ȉuĉU��M��U�H�E�H��H���������H�<I�߸    I�Ϟ������I�A��H�E�H��I��H�W�������H���H�E�H�E� �E�H�E� 9E�u��H��0[A_]���UH��AWSH�� ��H�����I��      L�H�}�H�u�H�E�� ��u�    �LH�E�� <wuH�E�H��I��H�a�������H���H�U�H�E�H��H��I��H�V.������H���H�E�H�E�H�� [A_]���UH��AWH����H�����I�i      L�H�}�H�U�H��I��H��/������H���H��A_]���UH��AWH����H�����I�      L�H�}�H�U�H��I��H��.������H���H��A_]���UH��AWH����H�����I��~      L؉}�H�u�H�M��U�H�Ή�I��H�0������H���H��A_]���UH��AWSH�� ��H�����I�~      L�H�}�H�}� u������VH�E�H��I��H�;2������H��ЉE�H�E؋@��u+H���������H�H��E�H�։�I��H�0������H��ЋE�H�� [A_]���UH��AWH����H�����I��}      L؉}�H�u�H�M��U�H�Ή�I��H��������H���H��A_]���UH��AWH����H�����I��}      L�H�}�H�U�H��I��H�r�������H���H��A_]���UH��AWSH��@��H�����I�I}      L�H�}ȉu�H�U�H�}� u	H�E��  H�E�H�E�H�E�H�E��E�    H�E�H��I��H�;2������H��ЉEԃ}����   H�E��@��u7�}�u�}� ~+H���������H�H��E�H�։�I��H�0������H��Ѓ}�
tk�E�;E�}E�}�u�}� ~H�E�H;E�vH�m��m��:�}��^���H�E�H�PH�U�UԈ�E��D����}�u�}� ~�m���E��)�������}�~	H�E��  ��Eԉ�H�E�H�E�H��@[A_]���UH��AWSH�� ��H�����I��{      L�H�}�H�u�H�}� u�    �^�E�    �2�E�Hc�H�E�H�� ��H�U�H�։�I��H��������H��ЃE�H�E�H��I��H�su������H��ЋU�9�w��E�H�� [A_]���UH��AWH��(��H�����I�K{      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I�
4������I�A��H��(A_]���UH��AWH��(��H�����I��z      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I��4������I�A��H��(A_]���UH��AWH����H�����I��z      L�H�}�H�U�H��I��H��Z������H���H��A_]���UH��AWH����H�����I�Fz      L�H�}�H�U�H��I��H��6������H��ҐH��A_]���UH��AWH��(��H�����I��y      L�H�}�H�u��U܋U�H�u�H�M�H��I��H�5������H���H��(A_]���UH��H����H�����I��y      L�H�}�H�}� u������!H�E��P#H�E���+  9�r�������    ����UH��AWH����H�����I�Hy      L�H�}�H�U�H��I��H�]6������H���H��A_]���UH��AWSH��`  ��H�����I��x      L�H������H������H�������E�    �E�    �  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H���������H���	E�}���  �E�H��    H��l  H�H��l  H�>��H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E��E�H������H�։�I��H�
�������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�}� t(H������H�E�H��H��I��H��������H����O  H������H��H���������H�<I��H��������H����   H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E�H�������E�H�։�I��H�Ȯ������H���H������H������H��H��I��H��������H����w  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������
   H��H��I��H�B�������H���H������H������H��H��I��H��������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������   H��H��I��H��������H���H������H������H��H��I��H��������H����  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�EȾ   H��fHn�I��H���������H���H������H������H��H��I��H��������H����]  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eк
   H��H��I��H���������H���H������H������H��H��I��H��������H����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ
   H��H��I��H�B�������H���H������H������H��H��I��H��������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ   H��H��I��H�B�������H���H������H������H��H��I��H��������H����G  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�E�   H��fHn�I��H���������H���H������H������H��H��I��H��������H����   H������H�ƿ%   I��H�
�������H��ЋE�Hc�H������H�� ��H������H�։�I��H�
�������H����4�E�Hc�H������H�� ��H������H�։�I��H�
�������H��ЃE��E�Hc�H������H�� ��������    H��`  [A_]���UH��H����H�����I�np      L؉��E��E�    �E��S��%wa��H��    H��e  H�H��e  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��o      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��H�� ��H�����I��n      L�H�}�H�u�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E�����UH��AWSH��  ��H�����I�gn      L�H������H������H��x����E�    H������H�E�f�E�  �E� �E�    �/  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H�\�������H���	E܃}���  �E�H��    H�Ed  H�H�:d  H�>��H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E��E�H�U�H�E�H��H��H��������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H�}� t'H�U�H�E�H��H��H��������H���H�E��e  H�E�H���������H�4H��H��������H���H�E��7  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E�H�������E�H�։�I��H�Ȯ������H���H������H�E�H��H��H��������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������
   H��H��I��H�B�������H���H������H�E�H��H��H��������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������   H��H��I��H��������H���H������H�E�H��H��H��������H���H�E��3  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�E��   H��fHn�I��H���������H���H������H�E�H��H��H��������H���H�E��x  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�E��
   H��H��I��H���������H���H������H�E�H��H��H��������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ
   H��H��I��H�B�������H���H������H�E�H��H��H��������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ   H��H��I��H�B�������H���H������H�E�H��H��H��������H���H�E��e  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�Eо   H��fHn�I��H���������H���H������H�E�H��H��H��������H���H�E��   H�E�H���������H�4H��H��������H���H�E�fǅ����  �E�Hc�H������H�� ������H������H�E�H��H��H��������H���H�E��8�E�Hc�H������H�� �E�H�U�H�E�H��H��H��������H���H�E��E��E�Hc�H������H�� �������H�E��  H�U�H������H)�H��H�Ā  [A_]���UH��H����H�����I��e      L؉��E��E�    �E��S��%wa��H��    H��\  H�H��\  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��d      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H���������L��Љ�<�����<���Hc�H�����H��  ��<���H���   A_]���UH��AWH���   ��L�����I��c      M�H����������H�����H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H����������H�����H��M��H���������L��Љ�<�����<���H���   A_]���UH��AWSH��0��H�����I��b      L�H�}؉u�H�U�H�M��}�   v
�    �   H�U�H�E�H��H��       H�<I��H���������H��ЉE�}���  ~�   �I�E�E�}� ~:�U�H�E�H��       H�4H��I��H��o������H��ЋE�Hc�H�E�H��  �E�H��0[A_]���UH��AWH����H�����I�%b      L؉}�H���������H�H�
�U�H�Ή�I��H��������H���H��A_]���UH��AWSH�� ��H�����I��a      L�H�}�H�}� tj�E�    �?H���������H�H��E�Hc�H�E�H�� ��H�։�I��H��������H��ЃE�H�E�H��I��H�su������H��ЋU�9�w���H�� [A_]���UH��AWH���   ��L�����I� a      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I�+`      M�H��8���H��0���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�H���������I�<M�׸    H�Ϟ������L�������UH��AWH����H�����I��_      L�H�}�H�U�H��I��H�)�������H��ҐH��A_]���UH��AWH��(��H�����I�A_      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H���������H��Ѹ    H��(A_]���UH��AWH��(��H�����I��^      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H���������H����H�E�H�E�� < tH�E�H   H9E�sH�E�� <
u�H�E��  H�E�H;E�����H��(A_]���UH��AWSH��0��H�����I�9^      L�H�}�H�uЉỦM�H��      H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H���������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H��      H�H�E�H��      �0H��      �D �}�u-�U�H�E�    H��I��H�w�������H���H�U�H��   �}�u+�U�H�E�    H��I��H���������H��Љ�H�EЉ�[�}�u,�U�H�E�    H��I��H���������H��Љ�H�E�f��)�U�H�E�    H��I��H���������H��Љ�H�EЈ�    H��0[A_]���UH��AWSH��0��H�����I��\      L�H�}�H�uЉỦM�H��     H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H���������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H��     H�H�E�H��     �0H��     �D �}�u'H�E�H��I��H���������H����Z�H�E�� �+�}�u%H�E�H��I��H���������H���fH~�H�U�H��    H��0[A_]���UH��SH��8��H�����I�Z[      L�H�}�H�u�H�U��E�    �E�    ��  �E�    �E�Hc�H�E�H�� ������%��  �E��E�Hc�H�E�H�� ������lu�E��E�   �E�Hc�H�E�H�� ����H���������H���	E�}��o  �E�H��    H�gS  H�H�\S  H�>��H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H���������H�����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H��������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�\�������H����?  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H�����   H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H����jH�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�\�������H������E��E�Hc�H�E�H�� ��������E�H��8[]���UH��H����H�����I��V      L؉��E��E�    �E��S��%wa��H��    H�VP  H�H�KP  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I�PV      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I�eU      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��H����H�����I�uT      L؉}�H�u�H�}� u������w�}��u������jH�E��@#��tH�E��@#�P�H�E��P#H�E��@#H�U��J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U���E�����UH��AWSH����H�����I��S      L�H���������H�H� H��I��H�;2������H��ЉE�}��t+H���������H�H��E�H�։�I��H�0������H��ЋE�H��[A_]���UH��AWH��(��H�����I�4S      L�H�}�H�u�H�U�H���������H�<I�ϸ    H�Ϟ������H�������UH��H����H�����I��R      L�H�}��	   H�E�H���r�����UH��SH����H�����I��R      L�H�}�H�}� u.H��     H�<H��������H���H��     H��H�E�H��H��������H���H�E�H��[]���UH��AWSH��0��H�����I�!R      L�H�}�H�u�H�E�H���������H�4H��I��H��������H���H�E�H�}� u
������   �E�    H�E�H��I��H�su������H��ЉE܃}�`~	�E�   �$H�E�H�P+H�E�H��H��I��H��r������H���H�E��@���H�E��PH�E�H��I��H���������H��ЋE�H��0[A_]���UH��H��0��H�����I�,Q      L؉}�H�u�H�E�H�E��E܉E��E�    �}� y,H�E�H�PH�U�� -�}�   �u�E�����E���E��؉E�H�E�H�E�M�Hc�Hi�gfffH�� ��������)�����)��ʉЍH0H�E�H�PH�U�ʈ�E�Hc�Hi�gfffH�� ����)ЉE�}� u��}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWSH��@��H�����I��O      L�H�}�H�u��U�H�}� u#H�E�H�E�H�E�H�PH�U�� 0H�E��  �  H�E�H�E؋E�Hc�H�E�H�H�E��3H�E؃��E�H�m��}�	~�7   ��0   �U��H�m���H�E�H�E�H;E�wËE�Hc�H�E�H��  H�E�H�E��E�    �8H�E�� <0uH�E��"H�U�H�E�H��H��I��H��r������H�����E��E�;E�|�H�E�H�E�H�E�H��I��H�su������H��Љ�H�E؋E�H�U�)Љ�H�M�H�E�HȾ    H��I��H�p������H���H��@[A_]���UH��AWH����H�����I�nN      L؉}�U�    ��I��H�y`������H���H��A_]���UH��AWH����H�����I�!N      L؉}�u�U��U��I��H���������H���H��A_]���UH��AWH����H�����I��M      L�H�}�H�U�H��I��H��c������H��ҐH��A_]���UH��AWH����H�����I��M      L�H�}�u�M�H�U��H��I��H��e������H���H��A_]���UH��H����H�����I�5M      L؉}�u�E��}�E��E��}�ЉE��}� x�E���y�E����E��E�+E�E��!�}� y�E���~�E����E��U��E�ЉE�H�E�����UH��H�� ��H�����I��L      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H�� ��H�����I�L      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H��H��H�����I�YK      L�H�}�H�u��U�H�E�H�E�H�E�H�PH�U�� ���E�E���H���������H�H������ ��uǃ}�-u�E�   H�E�H�PH�U�� ���E��"�E�    �}�+uH�E�H�PH�U�� ���E�}� t�}�u9�}�0u3H�E�� <xtH�E�� <XuH�E�H��� ���E�H�E��E�   �}� u�}�0u�   ��
   �E��}� t	H��   ������H�E�E�Hc�H�E�H�H��H�ЉE؋E�Hc�H�E�H�H��H�E�}� t�}� ~�E�)E�H�E��]�H�E�    �E�    �E���H���������H�H��������t�m�0�[�E���H���������H�H���������5  �E���H���������H�H��������t�7   ��W   )E�E�;E���   �}� ��   �}� tgH�E�H;E�|H�E�H;E�u0�E�;E�~(�E�����H�E�   �H���������H�� �����   �E�   �E�H�H�U�H��H�E��E�H�H)E��eH�E�H;E�H�E�H;E�u-�E�;E�~%�E�����H�E����H���������H�� �����$�E�   �E�H�H�U�H��H�E��E�H�HE���H�E�H�PH�U�� ���E��y������H�}� t�}� t
H�E�H���H�E�H�U�H�H�E�����UH��AWH����H�����I�%H      L�H�}�H�M�
   �    H��I��H���������H���H��A_]���UH��AWH����H�����I��G      L�H�}�H�M�
   �    H��I��H���������H���H��A_]���UH��AWAVAUATSH����H�����I�tG      L�H�}�H�uȉU�L�eп    L��L�`� �؉���H���������H�H������ ��uЃ�-u�   L��L�`� �����+uL��L�`� �؃}� t�}�u-��0u(A�$<xt	A�$<XuI�D$� ��I���E�   �}� u��0u�   ��
   �EċE�Hc������    H��I�ǋE�Hc������    H��H�Љ�A�    A�    ����H���������H�H��������t��0�T����H���������H�H��������tz����H���������H�H��������t�7   ��W   )�;]�}GE��x
M9�wM9�u��9�~A������A�   �E�H�L��Hc�I�L��L�`� ���;������E��yA�����H���������H�� "   �	����tI��H�}� tE��tI�D$��H�E�H�U�H�L��H��[A\A]A^A_]���UH��H����H�����I�1E      L؉}��   �   ���r����UH��AWSH����H�����I��D      L�H�}�H�E�H���������H�4H��I��H��q������H��Ѕ�uH���������H�H� ��    H��[A_]���UH��AUATSH�� ��H�����I�~D      L�H�}�H�u�H�8     ��E�L�e�H�]�E�,$L��L�`��H��H�XD�(�m��}� uې�H�� [A\A]]���UH��H��8��H�����I�D      L�H�}�H�u�H�U�H�8     ��E�H�E�H�E�H�E�H�E�H�E�H�E�H�E�� ���E�H�E�H�PH�U�H�U���H�E�H�PH�U�H�U���H�E�H�PH�U��U���m��}� u�������UH��SH��H��H�����I�YC      L�H�}�H�u�H�8     ��E�H�E�H+E��EȋE�9E���  �E�����EȺ    ��E��EȋU�H�E�H�H�E�H�E�H�E�H�E�H�E�E�H�H��H��H�E�H�H�E�H�E�H;E�sjH�0     H�H�U�H�E�H��H���щEă}� u/�E�H�H��HE�H�U�H�E�H��H��H�q�������H�����  �}� y�E�H�HE���  �H�E�H;E���   H�0     H�H�U�H�E�H��H���щEă}� u)�E�H�HE�H�U�H�E�H��H��H�q�������H���뢃}� ��   H�E�H;E�uA�E�H�HE�H�U�H�M�H�E�H��H��H��������H��ЋE�H�HE�H�E�H�E��M���H�U�H�E�H��H��H�q�������H��ЋE�H�H��HE��E�H�HE���   �E�H�H��HE�����H�E�H;E���   H�E�H+E�H��H�E�H+E�H9�|4�E�Hc�H�E�H�H�E�H��H��H���������H���H�E�H�E������H�U�H�E�H��H��H���������H��ЋE�Hc�H�E�H�H�E������E�H�H��HE�H�U�H�M�H�E�H��H��H��������H��ЋE�H�H��HE�H�E�H�E������H��H[]���UH��H�� ��H�����I�h@      L�H�}��u�U�H�M�H�0     H�U�H��U�H�8     ��U��U���H�U�H�H�U�H��H��H���������H��А����UH��AWH����H�����I��?      L�H�}�H���������H�<I�׸    H�Ϟ������H��Ѹ����H��A_]���UH��H��@��H�����I��?      L�H�}�H�u�H�U�H�U��H�E�H�U����H���������H�Hc���҃� ��u��E�    H�U���҃�+t��-u�E�   H�E�H� ���������E��E�    �E�    �E�    �;�M�H����������Y�H�U���҃�0�*��X��E�H�E��E�H�U����H���������H�Hc���҃���u�H�U����.uuH�E��?�M�H����������Y�H�U���҃�0�*��X��E�H�E��E��E�H�U����H���������H�Hc���҃���u��U�)U�}� uH� �������f���  �}� t�E�H��������f(fW��E�H�U����etH�U����E��   �E�    H�E�H�U���҃�+t��-u�E�   H�E��E�    �%�M܉����҉�H�U���҃�0ʉU�H�E�H�U����H���������H�Hc���҃���u��}� t�U�)U���U�U�}����|	�}�   ~H�����������   H����������E��E�E܃}� yF�]��A�E܃���t&�}� y�E��^E��E���E��YE��E��}��E��Y��E��}� u�H�}� tH�E�H�U�H��E�����UH��H����H�����I�V<      L؉}�H�E�   �E�    �H�U�H��H��H�H�H�E��E��E�;E�|�H�E�����UH��AWSH��@��H�����I��;      L��E�H�}��u�H�}� u	H�E��  H�E�H�E�H�(�������f��f/E�v,H�E�H�PH�U�� -�E�H�0�������f(fW��E��E�H�@�������f/s�E��H,�H�E��/�E�H�@���������\��H,�H�E�H�       �H1E�H�E�H�E�H�E�H��x�H*��H��H���H	��H*��X��M��\�f(��EȋE���H���������H���H��x�H*��H��H���H	��H*��X��YE�H�@�������f/s�H,�H�E��*H�@���������\��H,�H�E�H�       �H1E�H�E�H�E�H�M�H�U�H�E�H� �������H�43H��I�߸    I��������I�A��H�E�H��@[A_]���UH��AWH����H�����I�
:      L�H�}�H�U�    H��I��H�i�������H���H��A_]���UH��AWH����H�����I��9      L�H�}�H�u�H�M�H�U�H��H��I��H�i�������H����Z�H��A_]���UH��AWH��(��H�����I�`9      L�H�}�H�u�H�M�H�U�H��H��I��H�i�������H����E��E�H��(A_]���UH��H����H�����I�9      L؉}��E����3E�)�����UH��H��@��H�����I��8      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�    H�}� y>H�E�H�PH�U�� -H�       �H9E�uH��������H�E�H�E��H�E�H��H�E�H�E�H�E�H�M�H�gfffffffH��H��H��H��H��?H)�H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U��ʈH�M�H�gfffffffH��H��H��H��H��?H)�H��H�E�H�}� u�H�}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U߈H�E�H;E�w�H�E�����UH��AWH��8��H�����I�X7      L�H�}�H�uЉU�H�U�H�U�H�}� yH�U�H�JH�M��-H�]�H�U�H�U��}�u$H�M�H�u�   H��I��H��������H����H�M�H�U�H��H��H�$�������H���H�E�H��8A_]���UH��H��0��H�����I��6      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E�H�M�H���������H��H��H��H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U�ʈH�E�H���������H��H��H��H�E�H�}� u�H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWH��8��H�����I��5      L�H�}�H�uЉU�H�U�H�U�H�U�H�U��}�u$H�u�H�M�   H��I��H��������H����H�M�H�U�H��H��H�I�������H���H�E�H��8A_]���UH��H����H�����I�5      L؉}������UH����H�����I��4      Lظ   ]���UH��H����H�����I��4      L�H�}��    ����UH��H����H�����I��4      L�H�}�H���������H�H� ����UH��H����H�����I�b4      L�H�}�H���������H�H� ����UH��H�� ��H�����I�'4      L�H�}��u�H�U�H�M�    ����UH����H�����I��3      Lظ    ]���UH��H����H�����I��3      L��E�H�H�������f������UH��H����H�����I��3      L��E�H�H�������f������UH��H����H�����I�T3      L��E��}�H�H�������f������UH��H����H�����I�3      L��E�H�}�H�H�������f������UH��H����H�����I��2      L��E��M�H�H�������f������UH��H��(��H�����I��2      L��E��M��E��U��U��E��E��E������������������������������]��E�����UH��H����H�����I�/2      L��E����E����]��E�����UH��H����H�����I��1      L��E�H�P�������f������UH��H����H�����I��1      L��E�H�X�������f������UH��H����H�����I��1      L��E�H�`�������f������UH��H����H�����I�I1      L��E�H�h���������E��E�����UH��H����H�����I�1      L��E�H�p�������f������UH��H����H�����I��0      L��E�H�x�������f������UH��H����H�����I��0      L��E�H���������f������UH��H����H�����I�Z0      L��E�H���������f������UH��AWH����H�����I�0      L��E��E�H���������H�f(�fHn�I��H�W�������H���H��A_]���UH��H����H�����I��/      L؉}�H�u�    ����UH��AWH����H�����I��/      Lډ}�H�u�H���������H�<I�׸    H�Ϟ������H�������UH��AWH��(��H�����I�8/      Lى}�H�u�H�U�H���������H�<I�ϸ    H�Ϟ������H�������UH��AWSH�� ��H�����I��.      L�H�}�H���������H�<I�߸    H�Ϟ������H����E�    �.�E�H�H��    H�E�HЋ ��I��H�͝������H��ЃE��}�?~̸����H�� [A_]���UH��AWH����H�����I�E.      L�H�}�u�H���������H�<I�׸    H�Ϟ������H�����f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     �                                                                    ~ � � � � � � � � ~             ~ � � � � � � � � ~                 l � � � � | 8                   8 | � | 8                   < < � � �   <                < ~ � � ~   <                      < <              � � � � � � � � � � � � � � � �           < f B B f <           � � � � � � � � � � � � � � � �        2 x � � � � x             < f f f f <  ~               ? 3 ? 0 0 0 0 p � �              c  c c c c g � � �               � < � < �             � � � � � � � � � � �               > � >                  < ~    ~ <                f f f f f f f   f f              � � � {                | � ` 8 l � � l 8  � |                       � � � �              < ~    ~ <  ~              < ~                           ~ <                      �                         0 ` � ` 0                         � � � �                       ( l � l (                      8 8 | | � �                   � � | | 8 8                                                 < < <                  f f f $                             l l � l l l � l l           | � � � |   � � |               � �   0 ` � �             8 l l 8 v � � � � v           0 0 0 `                             0 0 0 0 0 0               0         0                   f < � < f                         ~                                    0                     �                                                           0 ` � �             8 l � � � � � � l 8              8 x       ~             | �    0 ` � � �             | �   <    � |               < l � �                 � � � � �    � |             8 ` � � � � � � � |             � �     0 0 0 0             | � � � | � � � � |             | � � � ~     x                                                       0                  0 ` 0                      ~     ~                     ` 0      0 `             | � �                       | � � � � � � � |              8 l � � � � � � �             � f f f | f f f f �             < f � � � � � � f <             � l f f f f f f l �             � f b h x h ` b f �             � f b h x h ` ` ` �             < f � � � � � � f :             � � � � � � � � � �             <         <                   � � � x             � f f l x x l f f �             � ` ` ` ` ` ` b f �             � � � � � � � � � �             � � � � � � � � � �             | � � � � � � � � |             � f f f | ` ` ` ` �             | � � � � � � � � |           � f f f | l f f f �             | � � ` 8   � � |             ~ ~ Z       <             � � � � � � � � � |             � � � � � � � l 8              � � � � � � � � � l             � � l | 8 8 | l � �             f f f f <     <             � � �   0 ` � � �             < 0 0 0 0 0 0 0 0 <               � � � p 8                 <         <          8 l �                                                   �       0                                     x  | � � � v             � ` ` x l f f f f |                   | � � � � � |                < l � � � � v                   | � � � � � |              6 2 0 x 0 0 0 0 x                   v � � � � � |  � x       � ` ` l v f f f f �                 8      <                        f f <       � ` ` f l x x l f �             8         <                   � � � � � � �                   � f f f f f f                   | � � � � � |                   � f f f f f | ` ` �             v � � � � � |                � v f ` ` ` �                   | � ` 8  � |              0 0 � 0 0 0 0 6                    � � � � � � v                   � � � � � l 8                   � � � � � � l                   � l 8 8 8 l �                   � � � � � � ~   �             � �  0 ` � �                 p                                        p         p                       v �                        8 l � � � �                               ��� ��� ~~~                                 uuu ��� ��� ���                                 ��� ��� ��� ��� ;;;                          ��� ��� ~~~ ��� ���                         ��� ��� ���     ��� ���                         ��� ���      ��� ��� ppp                 @@@ ��� ���         III ��� ���                 ��� ��� ��� ��� ��� ��� ��� ���                 ��� ���                 zzz ��� ���         ``` ��� ���                     ��� ���         ��� ��� MMM                     ��� ��� bbb     ��� ���                         ||| ��� ���      ��C@~Terminal shell.bin  BitMAP error
 Not suport BitMAP 4-bit Not suport BitMAP > 8-bit ____ none
 File name      KIB MiB GiB ./ File %s %lf            �@      �A      0AEntrada maior que o limite
 Erro ao criar o arquivo "%s"
       Error ao criar o arquivo "%s", atingio o limite de arquivos na entrada de directorio
   Panic: __malloc, sem espaco na tabela de alocacao
      panic: realoc sem espaco, %lx size = %d %d
 PWD strerrorr
      (((((�AAAAAABBBBBB                                �Dubug: %s %x %x
        (null)  ��������%���������������f����������������������m�������m�����������������������������������������������������������������������������������������������)�������ۗ��������������?�������?�������]���������������������������������������x���������������������������������������������������������������������������������������T�������f���������������������������������������f�������������������������������������������������������������������������������]���������������o�����������������������x�������(null) %        ��������̛������W����������������������h�������������������������������������������������������������������������������������������������������������џ��������������3���������������������3�������i�������i�������i�������i�������N�������i�������i�������i�������i�������i�������i�������i�������i�������i�������i�������*�������<�������i�������`�������W�������i�������<�������i�������i�������i�������i�������i�������i�������i�������i�������i�������3�������i�������E�������i�������i�������N�������panic: sscanf()
        �����������������������t����������������������L�������L�������������������������������������������������������������������������������������������������������$�������������������������������į��������������������������������������߯����������������������������������������������������������������������������������������������ͯ������������������������������������ͯ������������������������������������������������������������������������������į��������������֯����������������������߯������panic: freopen()
 r+ PWD call system funtion error. 
                 $@       �        %lu.%lu                �              �C                                                                        �_�
�@panic: signal()
 panic: sigaction()
 panic: setjmp()  panic: longjmp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �C �     �     �   �T �   �C �   �T �   �C �      �   �C �      �   �C �    4 �   �C �   D �                                   �2 �   �2 �   �2 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  zR x�  ,      @����   E�CG����B�A�          L   ����1   E�CG��     l   �����    E�C�� $   �   s���   E�CE��A�   $   �   `����    E�CG����B�A�$   �   �����    E�CG����B�A�(     �����   E�CG����B�A�   (   0  ���j   E�CG��W�B�A�       \  B����    E�CE���� (   �  ����   E�CG���B�A�       �  �����    E�CE���� (   �  e����   E�CG��q�B�A�   $   �  ����   E�CG����B�A�   $  ����9    E�Cp�     D  ����+    E�Cb�     d  �����    E�C��     �  -����   E�CE����   �  ����I    E�C@�     �  ����u    E�CE�f�A�(   �  I����   E�CG����B�A�   (     �����   E�CG����B�A�   $   D  �����    E�CG����B�A�,   l  j���2   E�CG���B�A�       (   �  l���D   E�CG��1�B�A�   $   �  �����    E�CG����B�A�(   �  �����   E�CG����B�A�   ,     ����   E�CG����B�A�       ,   L  a���   E�CG���B�A�       (   |  O����   E�CG��s�B�A�   $   �  �����    E�CG����B�A�(   �  h���   E�CG��
�B�A�   $   �  Y����    E�CG����B�A�$   $  ����   E�CF��A�   (   L  �����   E�CG����B�A�   $   x  G����    E�CG����B�A�(   �  ����5   E�CG��"�B�A�   $   �  ���k    E�CG��X�B�A�   �  K����    E�C��      �����    E�C��    4  ����X    E�CO� ,   T  ����l   E�CG��Y�B�A�       ,   �  ���6   E�CG��#�B�A�       (   �  ���D   E�CG��1�B�A�   (   �  %���q   E�CG��^�B�A�   (     j����   E�CG����B�A�   (   8  .���   E�CG����B�A�   (   d  ���Z   E�CG��G�B�A�      �  ���   E�C�   �  ����    E�C��    �  I���    E�C��     �  ���p    E�CF�`�A�$     ���    E�CG����B�A�$   <  ���r    E�CG��_�B�A�(   d  '��   E�CG��	�B�A�   $   �  
���   E�CF���A�       �  ����    E�CE���A�    �  [���    E�CE���A�    	  ����    E�C��     	  ���A    E�Cx�      @	  ���i    E�C`�        d	  ��U    E�CL�    �	  D��U    E�CL�    �	  y��i    E�C`�    �	  ���g    E�C^�    �	  	���    E�C�� $   
  ����   E�CE�{�A�      ,
  2��9    E�Cp�  $   L
  K���    E�CG����B�A�   t
  ��^    E�CU� (   �
  J��   E�CG���B�A�   (   �
  3���   E�CG����B�A�   (   �
  ���]   E�CG��J�B�A�   (     ��   E�CG��l�B�A�   (   D  U��D   E�CJ��.�B�A�   (   p  m"��:   E�CG��'�B�A�   $   �  {#��    E�CG����B�A�   �  S$���    E�C��    �  %���    E�C�� (     �%���   E�CJ����B�A�   (   0  ~)��i   E�CG��V�B�A�   (   \  �,��H   E�CG��5�B�A�   (   �  �.��e   E�CJ��O�B�A�      �  3��a    E�CX�    �  Q3��9    E�Cp�      �  j3���    E�CF�w�A�(     �3��'   E�CG���B�A�   $   D  �6��   E�CE���A�   $   l  �8���   E�CF���A�      �  :��    E�C��    �  �:���    E�C�� (   �  �;��O   E�CG��<�B�A�   $      �<���    E�CG����B�A�(   (  �=��C   E�CG��0�B�A�      T  �?��k    E�Cb� $   t  @���    E�CG����B�A�   �  �@���    E�C��    �  >A��w    E�Cn�    �  �A��b    E�CY� $   �  �A���    E�CG����B�A�$   $  jB��z    E�CG��g�B�A�   L  �B��a    E�CX�    l  �B���    E�C��    �  wC��{    E�Cr� $   �  �C��+   E�CF��A�      �  �D��6   E�C-�   �  �E��L    E�CC� $     F���    E�CG����B�A�   <  �F���    E�Cw�    \  G��}    E�Ct� $   |  tG��r    E�CF�b�A�    $   �  �G���    E�CF���A�       �  )H���    E�C��    �  �H��3   E�C*�     �I��7   E�C.�   ,  �J��W    E�CN� $   L  'K���    E�CG����B�A�$   t  �K���    E�CG����B�A�   �  L���    E�C�� $   �  �L��V    E�CF�F�A�       �  �L��P    E�CF�         M��U    E�CL�    $  DM��U    E�CL� $   D  yM���    E�CG����B�A�$   l  �M���    E�CG����B�A�$   �  aN��K    E�CF�{�A�     $   �  �N��K    E�CF�{�A�     $   �  �N��S    E�CF�C�A�    $     �N���    E�CG����B�A�$   4  BO��S    E�CF�C�A�    $   \  mO��K    E�CF�{�A�     ,   �  �O��[   E�CG��H�B�A�       $   �  �P���    E�CG����B�A�$   �  7Q��]    E�CF�M�A�    $     lQ��]    E�CF�M�A�    $   ,  �Q��K    E�CF�{�A�     $   T  �Q��L    E�CF�|�A�     $   |  �Q��Y    E�CF�I�A�       �  R��Y    E�CP� $   �  RR��K    E�CF�{�A�     (   �  uR���   E�CJ��{�B�A�         �Z���    E�C��     $   <  `[���    E�CI���A�       d  #\��l    E�Cc� (   �  o\���   E�CJ����B�A�       �  e���    E�C��     $   �  �e��   E�CI���A�    $   �  wf���    E�CI���A�    $   $  <g���    E�CG����B�A�$   L  �g��\    E�CF�L�A�    $   t  !h���    E�CG����B�A�$   �  �h���    E�CI���A�       �  li���    E�CI�    $   �  �i��L    E�CF�|�A�           j��e    E�CF�U�A�    0  Rj���    E�CF���A�(   T  �j���   E�CG����B�A�   (   �  Hl��=   E�CG��*�B�A�   $   �  Ym��\   E�CE�M�A�      �  �q���    E�C�� $   �  r���    E�CI���A�    $     �r���    E�CI���A�       D  �s���    E�C�� $   d  9t���    E�CG��z�B�A�   �  �t��Y    E�CF�       �  �t��9    E�Cp�  $   �  �t���    E�CE�q�A�    $   �  Hu���    E�CG����B�A�     v��G   E�C>�,   <  ?w��u   E�CG��b�B�A�       $   l  �x��M    E�CF�}�A�     $   �  �x��O    E�CF��A�     $   �  �x��L    E�CF�|�A�     $   �  �x��S    E�CF�C�A�         y���    E�C�    ,  �y���    E�C��    L  z���    E�C��    l  �z��2   E�C)�$   �  �}��U    E�CF�E�A�    $   �  �}��U    E�CF�E�A�    4   �  ~��L   E�CM�����-�B�B�B�B�A�        ���7    E�C       $   4  2���w    E�CG��d�B�A�(   \  ����{    E�CI���d�B�B�A�   �  Ѐ���    E�C�� $   �  ^����   E�CE���A�       �  (����    E�Cx�     $   �  ����\    E�CF�L�A�         ����5   E�C,�   <  ·��_    E�CV� ,   \  ����   E�CG����B�A�       $   �  ȉ��P    E�CF�@�A�    $   �  ����Z    E�CF�J�A�    $   �  "���^    E�CF�N�A�         X���4    E�Ck�     $  l���v   E�Cm�$   D  ���    E�CF���A�       l  I����    E�C�� $   �  "����    E�CF���A�       �  ����*    E�Ca�     �  ����'    E�C^�     �  ����/    E�Cf�       ����;    E�Cr�     4  ʍ��;    E�Cr�     T  ���:    E�Cq�     t  ����'    E�C^�     �  ���9    E�Cp�     �  ���9    E�Cp�     �  8���<    E�Cs�     �  T���=    E�Ct�       q���>    E�Cu�     4  ����n    E�Ce�    T  ݎ��;    E�Cr�     t  ����9    E�Cp�     �  ���9    E�Cp�     �  *���9    E�Cp�     �  C���D    E�C{�     �  g���9    E�Cp�        ����9    E�Cp�     4   ����9    E�Cp�     T   ����9    E�Cp�  $   t   ˏ��a    E�CF�Q�A�       �   ���2    E�Ci�     �   ���T    E�CF�   �   N���X    E�CF�$   �   �����    E�CG����B�A�   !  ����T    E�CF�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            GCC: (Ubuntu 9.3.0-17ubuntu1~20.04) 9.3.0                                        �                    �                  @ �                 p@ �                 �@ �                 �@ �                  ` �                                     ��                     ��_ cole _             ��                )        �           P         �           0    ��                7    ��                >      h2 �           C      s2 �           H    ��                N    ��                Y    ��                b    ��                >      ~2 �           C      �2 �           h      �2 �           m    ��                t    ��                }    ��                �     �E  �         �    ��                �    ��                >      �2 �           �    ��                �     �@ �          |    �@ �          �     �@ �          >      �2 �           �    ��                �    ��                >      �2 �           �    ��                �    ��                �     �@ �           �      A �           �     �@ �          �     ze  �   �      �     jh  �   �           �2 �           	     �2 �                �2 �                �2 �                 3 �                3 �           "     �2 �           '     �2 �           -   ��                4   ��                >      3 �           C      ,3 �           h      P3 �           �   ��                :     A �          >      �3 �           C      �3 �           J   ��                Q   ��                >      4 �           X   ��                a   ��                j   ��                s   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                   ��                    (A �             ��                $   ��                -   ��                7   ��                A   ��                >      4 �           L   ��                T   ��                ^   ��                h   ��                >       5 �           p   ��                x   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �    ��  �   �       >      85 �           �   ��                �   ��                �    ��  �   �       >      07 �           C      77 �           �   ��                �   ��                �   ��                	    @A �             ��                �   ��                �   ��                   ��                >      09 �           #   ��                ,   ��                6    !�  �   e       h    ��  �   �       K    (�  �   �      @    @A �          J    ��  �   =      Q    @B �          �    e�  �   �       -   ��                .   ��                [   ��                d   ��                n   ��                >      8; �           x   ��                �    @C �   `       �   ��                >      J; �           �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                >      M; �           �   ��                    �C �              �C �              ��  �   {           \�  �   �           
�  �   �      !   ��                >      Q; �           *   ��                >      p; �           C      x; �           h      �; �           3   ��                :     �   _       >      �; �           C      �; �           h      �; �                �; �           E   ��                L   ��                U   ��                _   ��                e   ��                l   ��                s   ��                t   ��                {   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                >      �; �           �   ��                �   ��                �   ��                >      �; �           �   ��                >      �; �           �   ��                >      �; �           �   ��                >      �; �           �   ��                >      �; �           �   ��                >      �; �           �   ��                >      �; �           �   ��                >      �; �           �   ��                >       < �           �   ��                �   ��                >      < �           C      < �           �   ��                >      -< �           C      >< �                ��                    p@ �                �   T       "    �|  �         �    =�  �   \       5    <L  �         ?    �)  �   �       J    �  �   {       Q    � �   9       U    5 �   ;       Z    � �   �       a    �{  �   �       q    �;  �   �       u    �  �   7      L    ?�  �   �       ~    �C �          �    ��  �   �      �    ��  �   �       �      �               %  �   �       �      �           �    Ǿ  �   P       �    �	 �   �       �    �T �          �    ��  �   �       �    w�  �   �       �    �C �          �    �  �   �      �    ��  �   U       �    �5  �   u       �    j�  �   w       �    
 �   9       �    �T �          �    � �   9       �     �   ^           `2 �              ��  �   �       =    �  �   �           �  �   [          �  �   :      &    �  �   �       6    	d  �   q      v
    ��  �   �       B    ��  �   w       �    �I  �   �      I    (2  �   �       X    9  �   �      `    ��  �   L       g    � �   v      �    ��  �   �       n    �  �   U       v    }  �   \       }    ��  �   Y       �    ��  �   M       �    ��  �   K       
    �C �          �    `L �          �    Z  �   �       �    �2  �   �      �     �   <       �    d�  �   �       �    �B  �   �      �    ��  �   L      �    8�  �   G      �    �C �          �    Wl  �         �    ��  �   ]          �%  �   �       8     L �   4           D�  �   K              �               �&  �   �      $    96  �   �      +     ` �           4    �j  �   Z      >    �  �   �       D    �v  �   A       K    /�  �   �       W    �<  �   2      ^    �^  �   6      e    ;u  �   �       m    �  �   2      t    �C �          y    @�  �   �       �    6o  �   �       �    f�  �   �       �    PB  �   �       �    �
 �   �       �    A�  �   O       �    �  �   5      �    �G  �         �    w  �   i       �    #[  �   l      �    X �   P       K    ��  �   �       �    �W  �   5      �    �u  �   �       �    ��  �   z       �    �~  �   �      a     � �                ��  �   �           h�  �   Y           Q  �             )�  �   9       ,    Ñ  �   �      5    m �   �      )    � �   9       :    �C �          @       �          k
    �@ �           I    �T �          O       �           V    �C �          _     � �           e    w�  �   �       l    b{  �   9       v    �x  �   g       �
     �   D       �	    q �   '       �    � �   >       �    � �   T       �    q�  �   V       �    ��  �   �       �    �w  �   U       �    $  �         �    � �   n       �    w�  �   }       �    m#  �   �       �    װ  �   �       �    � �   9       �    �L �          �    ��  �   S       �    8(  �   j      	    �  �   k       	    �  �         l
    �@ �           	     �  �   W        	    �  �   H      +	    h�  �   �       2	    4�  �   �       9	    ��  �   �       E	    �  �          P	    ��  �          [	    * �   X       e	    zt  �   �       l	    �  �   �       �    @  �   D      }	    �  �   ]       �	     4 �          �	    ��  �   D      �	    �T �          �	    �y  �   �      �	    �  �   �       �	    c�  �   �       
       �           �	    ��  �   9       �	     �   ;       �	    u�  �   b       �	    �C �          �	    <"  �   1      �	    �  �   K       �	    G �   *       �	    YP  �   �       �	    ��  �   K       �	    ��  �   �           � �   /       
    p  �   r       
       �           
    �C �          �    ��  �   �       �    C �   a       
    �  �         �
    ��  �   S       (
    �1  �   +       �    �r  �   �      6
    n  �   �       >
    ��  �   l       7    �p  �         H
    m�  �   �       q
    _ �   9       O
    {5  �   I       U
    �Z  �   X       ^
    c�  �   e      j
    �@ �           p
    p �   9       u
    ��  �   K       �    v�  �         {
    ^*  �         �
    � �   Z       �
    ��  �   6      �
    � �   9       �
    
	 �   �       �
    � �   2       >    ��  �   �       �
    �C �          �
    ��  �   i      �
    ��  �   �       �
    um  �   �       �
    �  �   '          ��  �   �       
       �           �     D �          �
    z�  �   S       �
    �n  �   p       �
     0 �   @      �
    N   �           �
    ҫ  �   C          = �   :           �  �   u          a�  �   �           t�  �   ]            "R  �   �      ,    D �          `     � �           5    �X  �   k       <    	�  �   \      D    �  �   L       K    .�  �   Y       S    CY  �   �       �       �           ]    ��  �   �       g    3�  �   7       l    D �          s    �V  �   �       �    ȟ  �   a       �    =�  �   U           �0  �         �    b�  �   �       �     D �          .    9,  �   �      �    !x  �   i       �    � �   ;       �    ��  �   3      �    `   �   �      �    }+  �   �       �    �  �   L       �       �           �    l�  �   U       �    �1  �   9       �    �x  �   �       �    UK  �   �            w �   '       �       �               �|  �   ^           /�  �   �           ` �   4           �  �   a       "    s�  �   �       (    � �   9       -    ��  �   +      7    �a  �   D      D    L �   =       J    e�  �   �      S    ��  �   r       [    ww  �   U       g    ��  �   L       l    ��  �   O       lib/setup.asm HEADER_MAGIC HEADER_FLAGS header crt0.c term.c .LC0 .LC1 gui.c font8x16.c window.c bmp.c .LC2 font.c border.c editbox.c editbox_refresh mouse.c menubox.c obj.c objm foc message.c dialog.c button.c listbox.c file_data file_type file_unidade attr .LC3 .LC4 .LC5 .LC6 .LC7 .LC8 .LC9 .LC10 file.c cfs.c alloc_spin_lock pipe.c path.c memcmp.c memcpy.c memset.c strcasecmp.c strcat.c strchr.c strcmp.c strcpy.c strcspn.c string.c strlen.c strncasecmp.c strncmp.c strncpy.c strpbrk.c strrchr.c strsep.c strspn.c strtok.c last.1481 strstr.c strdup.c memmove.c strcoll.c strerror.c ctype.c tolower.c toupper.c stdio.c fopen.c fclose.c fflush.c fputc.c fgetc.c fgets.c fputs.c fread.c fwrite.c remove.c rewind.c fseek.c feof.c ftell.c vfprintf.c vf vsprintf.c vsnprintf.c sn_buf putchar.c sscanf.c perror.c vfscanf.c character _buf.1638 fvalue _buf.1650 ungetc.c getchar.c freopen.c tmpnam.c _tmpnam rename.c itoa.c i2hex.c malloc.c calloc.c free.c realloc.c lldiv.c strtol.c atoi.c atol.c strtoul.c exit.c getenv.c qsort.c qscmp qses qsexc qstexc qs1 system.c strtod.c ftoa.c _precision atof.c strtof.c strtold.c abs.c ltoa.c utoa.c srand.c errno.c gmtime.c localtime.c strftime.c clock.c math.c pow.c sqrt.c atan.c acos.c asin.c floor.c ceil.c exp.c locale.c signal.c setjmp.c _GLOBAL_OFFSET_TABLE_ longjmp read_directory_blk menumotor drawstring strcpy log sqrt setjmp clean_blk_enter put strtok_r stdout vsprintf ungetc pwd_ptr argv strerror utoa_r __m_i memmove __tm __realloc_r atol __window_puts getenv ceil errno floor strtold _infinity qsort fgets file_update file_read_block m_file_list memcpy __window_clear BitMAP2 perror ltoa_r tolower system feof malloc remove fs_directory msg_read __window_putchar ldexp vsnprintf m_edit strtoul itoa __pipe__ stdgetc_r update_directory_entry _drawline fflush argc drawrect BitMAP eh_frame stdputc_r upath tell_r strncasecmp border button write_r strtol user rename flush_r strrchr update_editbox utoa calloc strtod fmouse rewind_r dialogbox atof update_objs seek_r strcat read_directory_entry debug_o fseek obj_focprocess __free_block_r open_dir ftoa stdin font8x16 __m_c _start obj_list __end strstr write_blk get_file_name atan2 signal strcoll strncmp write_sector draw_char_transparent pow strncpy put_pixel strcasecmp log10 _BLK_ realloc drawchar path_count open_file_r strtok remove_blk memcmp sscanf getfilename file_close pipe_write sigaction read_r file_write_block fread _ctype open_file addr search_blk_null strdup fopen sysgettmpnam localtime memset pwd main ftell srand init_process fclose getchar close_r __data ptr_mouse2 __free_r update_window getkeyw _vsputs_r strcmp color msg_init remove_file __bss atan fgetc drawchar_trans strtof strcspn asin ltoa setlocale stderr create_file strsep getkey __malloc_r fputc open_r A__ call_function getpathname strftime i2hex lldiv fwrite obj_process __window getmsg vfscanf rewind freopen msg_write pipe_read exit pipe_r register_obj __block_r atoi __heap_r ptr_obj assert_fn gmtime strspn ctr0 drawstring_trans strlen __code toupper wcl filename_cmp submenubox clock read_super_block abs strchr fputs acos strchrnul file_listbox frexp vfprintf strpbrk read_sector free setpath  .symtab .strtab .shstrtab .text .data .got .got.plt .data.rel.local .bss .eh_frame .comment                                                                                        �                                       !                �                                          '              @ �    @     p                              ,             p@ �   p@                                  5             �@ �   �@                                   E             �@ �   �@     @                             J              ` �    P      0                             T      0                �     *                                                   0�     `-      
   �                 	                      ��     t                                                   �     ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ELF          >       �   @       ��         @ 8  @                   �      �    �       �                             �      �   0"       0                   0      0 �    0 �    0       0             Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��  ���_ cole _          �      �            ` �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           I��H�0% �   L�H�% �   H�H�   �   L�H�  �   L�#H�  �   L�+�   �����H��H��H��H��L�������UH��AWSH��@��H�����I���      L�H�}�H�u�H�U�H�M�L�E�L�M�H���������H�H�U�H�H��     H�E�H�H�E�H��     H�H��     H�H� H��H��     H�H��     H�H��H�x     H�H��     H�H�@H��H�p     H�H�E�H��     H�H�E�H�h     H�H�E�H��     H�H��     H�H��H��     H�I�߸    H�-f������H���H��     H�    H���������H�H� H��H��     H�H���������H�H� H��H���������H�H� H�։�I��H��������H��ЉE�E��I��H���������H��АH��@[A_]���UH����H�����I�$�      Lڸ    H��������H�
�Ҹ    ]���UH��AWSH����H�����I���      L�H�E�   �    H��I��H�@v������H���H���������H�H�H�E�H��H��I��H�~n������H����E�f=t�ǐ�H��[A_]���UH��AWSH��0��H�����I�S�      Lۉ}�H�u��}� 
������D  H�E�H� H�E�H�E�H�E�� <0u
������  H��     H�H�E�H�E�!  �    H��I��H�@v������H��ЋE�Hc�H�E�H�H�E�H�E�   �E�    �?�E�H�H��    H�E�H�H�H�E�H��H��I��H��x������H���H�E�   �E��E�;E�|�H��     H�H�U�H��H��I��H��x������H���H��     H�<H��     H�4H���������H�H� �   �   I���r�    H�������H��Ҹ    H��0[A_]���UH��H����H�����I���      L�H�}��E�    H�U�H�U��w�U��J�M�H�M�H��     Hc�H�H���H�E�H�U����tH�U���� u�H�U����t5H�U�H�JH�M�� �H�E�H�U���� t�H�U����t�}�~������E�����UH��AWSH�� ��H�����I��      L��E�    �   I��H���������H���H�E�   I��H���������H���H�Eؿ�   I��H���������H���H��     H��!  I��H���������H���H��H��     H��   �    H��     H�<I��H�@v������H���H�E�   �    H��I��H�@v������H���H�z�������H�<I��H�5�������H���H��H�E�H�~�������H�4H��I�߸    H�A�������H��ѿ �  I��H�7&������H���H�E�H��H���������H�<I�߸    H�
�������H��ҿ����I��H�7&������H���H���������H�H�H�E�   H��I��H��������H���H�E�H��H�)������H��ЉE�H��     H�H�E��E�    �]  H�}� �N  H�       �E�Hc�H�H��H�H�H��H�H�H�E�H��H��I��H�8x������H��Ѕ�ucH�       �E�Hc�H��H�H�H��H�H�H��H� H��H��     H�H��     H��E�H��     H�4�����   �}�u.H�E�H��H���������H�<I�߸    H�
�������H����qH�Eк   H���������H�4H��I��H��|������H��Ѕ�uAH��     H��������H�H�H��     H��E�H��     H�4������E��}�������7�����UH��AWH����H�����I���      L؉}�H�u�H���������H�<I��H�d�������H��Ҹ    H��A_]���UH��AWH����H�����I�4�      L؉}�H�u�H���������H�<I��H�d�������H��Ҹ    H��A_]���UH��H����H�����I���      L؉}�H�u�   �   ���r�    ����UH��AWSH����H�����I���      Lۉ}�H�u��}�~9H�E�H��H�H�E�H��H� H��H��I��H��������H��Ѕ�u�    �*H���������H�<I�߸    H�
�������H��Ҹ����H��[A_]���UH��H����H�����I���      L؉}�H�u�   �   ���r�    ����UH��AWSH�� ��H�����I���      Lۉ}�H�uЃ}�������^H�E�H��H� H���������H�4H��I��H�.�������H���H�E�H�}� u������H�E�H��I��H�Ć������H��и    H�� [A_]���UH��AWH����H�����I��      L؉}�H�u�H���������H�<I��H�d�������H��Ҹ    H��A_]���UH��AWSH��   ��H�����I���      Lۉ�l���H��`���H��p�����   �    H��I��H�@v������H���H��p���H��H���������H�<I�߸    H�
�������H��Ҹ    H�Đ   [A_]���UH��AWSH�� ��H�����I� �      Lۉ}�H�u�H��������H�<I��H�d�������H����E�    ��   H�       �E�Hc�H�H��H�H�H��H�H� H��I��H�d�������H���H�       �E�Hc�H�H��H�H�H��H�H� H��I��H��{������H��ЉE���    I��H��������H��ЃE��}�~�H�       �E�Hc�H�H��H�H�H��H�H��H� H��I��H�d�������H��п
   I��H��������H��ЃE��}�� ����    H�� [A_]���UH��H����H�����I���      L؉}�H�u�    ����UH��AWH����H�����I���      L؉}�H�u�H���������H�<I��H�d�������H��Ҹ    H��A_]���UH��AWH����H�����I�-�      Lډ}�H�u�I�׸    H�������H��Ѹ    H��A_]���UH��AWSH����H�����I���      Lۉ}�H�u��}�,H��������H�<I�߸    H�
�������H��Ҹ�����UH�E�H��H� H��I��H���������H��Ѕ�t,H��������H�<I�߸    H�
�������H��Ҹ������    H��[A_]���UH��AWH����H�����I��      L؉}�H�u�H���������H�<I��H�d�������H��Ҹ    H��A_]���UH��AWH����H�����I���      L؉}�H�u�H���������H�<I��H�d�������H��Ҹ    H��A_]���UH��AWH��(��H�����I�j�      L؉}�H�u�H���������H�H�H�U�H�U�H��I��H��"������H��Ҹ    H��(A_]���UH��AWSH��0��H�����I��      Lۉ}�H�u��}�
�    ��  H�E�H��H� H�<�������H�4H��I��H�8x������H��Ѕ�u!I�߸    H��p������H��Ҹ    �  �    I��H���������H���H�E�H�E�    �    H��I��H�@v������H��п   I��H���������H���H�E�H�E�H��H�H�E�H�?�������H�4H��I�߸    H�A�������H���H�M�H�E�@   H��H��I��H��W������H��ЉE�H�E�H��I��H�[�������H���H�E�H��I��H�[�������H��Ѓ}��u:H�E�H��H� H��H�H�������H�<I�߸    H�
�������H��Ҹ�����cH�E�H��H� H��I��H�bo������H��Ѕ�t:H�E�H��H� H��H�H�������H�<I�߸    H�
�������H��Ҹ������    H��0[A_]���UH��AWSH����H�����I���      Lۿ    I��H���������H���H�E�H�E�    �    H��I��H�@v������H���H�E�@   H��H�k�������H�<I��H��W������H��ЉE��}��uHH�n�������H�<I�߸    H�
�������H���H�E�H��I��H�[�������H��и    �'  �}� uHH�z�������H�<I�߸    H�
�������H���H�E�H��I��H�[�������H��и    ��   �E�    �   H�E��@b����@��t\� �� I��H�7&������H���H�E�H��H���������H�<I�߸    H�
�������H��ҿ����I��H�7&������H����,H�E�H��H���������H�<I�߸    H�
�������H���H�m考E��E�;E��Q���H�E�H��I��H�[�������H��и    H��[A_]���UH��H��0��H�����I���      L�H�}�H�u��U܉M�L�E�H���������H�H� H�E��E�H9E�}?H�E��@��H9E�}0H�E�H�E��E�H�E�H��H�E�H�H��    H�E�HE؉������UH��SH��@��H�����I�4�      Lۉ}ԉuЉỦM�L�E�L�M�f�E�  H�E�H�@H�E�H�E��@�E�}�u�E�    �E�    �   f�E� H�E��@�EȉE��H�H� H�E�H�� f�E�H�E�� ���E��J�E�f#E�f��t5�UЋE��Hc��UԋE��H�H�}��M�U�I��H��H�)������H���f�e�m��}� y��E�H�E��@9E��b�����H��@[]���UH��AWSH��0��H�����I��      Lۉ}܉u؉UԉM�D�E�L�M��E�    �X�E�    �CH�E�L��   �M�H�E��P�u؋E��Hc��}܋E��H�H��I��H�)������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I�n�      Lۉ}܉u؉UԉM�D�E�L�M��E�    �p�E�    �[H�E�H��   �E��E�i��E��A��H�E��P�M؋E��Hc��M܋E��H�I��D��H��I��H�)������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I���      Lۉ}܉u؉UԉM�D�E�L�M��}� �[  �}� �Q  �E�    �>H�E�L��   �M�H�E��P�E�Hc��}܋E��H�H��I��H�)������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E����Hc��}܋E��H�H��I��H�)������H��ЃE��E�;E�|��E�    �AH�E�H��   �M�H�E��P�u؋E��Hc��E�H�I��H��I��H�)������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E��Hc��}܋E����H�H��I��H�)������H��ЃE��E�;E�|���H��0[A_]���UH��AWSH��@��H�����I���      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}��  �E�    ��   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��   �E�f#E�f��tDH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�)������H����BH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�)������H���f�e�m��}� �[����E�H�E��@9E��	�����H��@[A_]���UH��SH��8��H�����I���      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H��������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I���      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}���   �E�    �   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��W�E�f#E�f��tBH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�)������H���f�e�m��}� y��E�H�E��@9E��T�����H��@[A_]���UH��SH��8��H�����I���      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H�������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I���      L�H�}ȉuĉU��M�D�E�D�M�H���������H�H� H�E�H�E�H   � �? �    H��I��H�@v������H����E�    �U�H�E��P4�UH�E��P8�UH�E��P<H�E��@H   H�E��@L   H�E��P<H�E��PP�UH�E��PTH���������H�H��H�E�H�PXH�E��@D    H�E��PDH�E��P@�U�H�E��P�U�H�E��P�U�H�E��P �U�H�E��P�U H�E��P`�} u�E�   H�E��@�P�H�E��P(H�E��P�E�)ЍP�H�E��P$H�E��@0   �E����H�E��P,H�E��@��H�E��@��H�E�I���Ѻ    �    I��H��-������H���H�E��@4��H�E��@����H�E�I��A�ȹ   �   �   H��������H��Ѓ}� u:H�E��@����H�E�I��A���� �   �   �   H��������H����8H�E��@����H�E�I��A���� �   �   �   H��������H��Ѓ}� t}H�E��@����H�U��E�I��A���� ����   �   H��������H���H�E��@4��H�E��@���ƋE��H�U�I��A�ȹ   ��ƿ   H��������H���H�E��@8A��H�E��@$��H�E��@(��H�E��@,��H�E��@0��H�E�I��H��������H���H�E�H��I��H��{������H������E�H�E�H�pHH�E��@��E܉������)Љ�H�E�H���u�I��A���� ������   ��H��H�9������H���H��H�E��@����H�E�I��A�    �   �   �   H�J������H���H�E�H�PHH�E��@��H���u�I��A���� ������   �ƿX   H�������H���H��H�E�H�PHH�E��@��(H���u�I��A���� ������   �ƿ-   H�������H���H��H�E�H�e�[A_]���UH��AWSH��0��H�����I�x�      L�H�}�H�u�H�E��P0H�E��@Ѓ�P�E�H�E��P,H�E��@Ѓ��E��E�P   �E�   �E�    �E���� H�E�H��I��H��{������H��ЉE�H�E�L�@H�M؋U܋E���������p��E�<�E��������ƋE���)ƋE��H�E�H���u�M��A�ȉщ�H��H�^������H���H���H�e�[A_]���UH��H����H�����I�t�      L�H�}��   H�E�H���r�����UH��H����H�����I�;�      L�H�}������UH��H����H�����I��      L�H�}�H�U��BD    H�U��JDH�U��J@H�U��R8A��H�U��R$��H�U��R(A��H�U��R,��H�U��R0��H�U�I��D��I��������J��А����UH��SH��(��L�����I���      Mډ�f�E�H���������I�H� H�E�H���������I�H��H�E�H�PXH�E�@(�P�H�E�@H���к    ��E�H�E�@$�P�H�E�@L���к    ��E�H�E�P<H�E�PPH�E�PD�E�9�rH�E��@D    H�E�@@�PH�E�P@H�E�P@�E�9�r9H�E��@D    H�E�PDH�E�P@H�E�H��H��"������I����E��  f�}���   H�E�@D����   H�E�@D�P�H�E�PDH�E�H�xHH�E�pTH�E�@PH�U�J,H�U�RLA��H�U�R@A��ʃ���H�U�J0H�U�RHA��H�U�RDA��ʃ�A��H���u�I��A������D�޿    H��������I���H����   f�}�	uH�E�@D�PH�E�PD��   f�}�
u!H�E��@D    H�E�@@�PH�E�P@�   f�}���   H�E�H�xHH�E�pTH�E�PPH�E�H,H�E�@LA��H�E�@@A��ȃ���H�E�H0H�E�@HA��H�E�@DA��ȃ�A���E�H���u�I��A���щ�D�މ�H��������I���H��H�E�@D�PH�E�PD�E�H�]�����UH��H����H�����I���      L؉}�H���������H�H� H�E��U�H�E��P<�����UH��SH��(��H�����I�s�      L�H�}�H�}� t=H�E�H�E��&H�E�H�PH�U�� f�����H�q#������H���H�E�� ��u���H��([]���UH��AWSH��P��H�����I���      L�H�}��u��U��M�L�E�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H���������H�<I�߸    H�
�������H��Ҹ�����6  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H���������H�<I�߸    H�
�������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H���������H�<I�߸    H�
�������H��Ҹ   ��   �E�    �   �E�    �   �}� tNH�E�H��   H�E��P�M��E���E��Hc��M��E���E��H��M�I��H��I��H�)������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�)������H��ЃE��}� �U����E��}� �;����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��P��H�����I��      L�H�}��u��U��M�D�E�L�M�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H���������H�<I�߸    H�
�������H��Ҹ�����3  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H���������H�<I�߸    H�
�������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H���������H�<I�߸    H�
�������H��Ҹ   ��   �E�    �   �E�    �   �}� tKH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�)������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�)������H��ЃE��}� �X����E��}� �>����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��0��H�����I�7�      Lۉ}܉u؉U�H�M��E�    �   �E�    �t�U�������E��H���������H�Hڋ��E�}� tBH�E�H��   H�EȋP�MԋE��Hc��M؋E��H��M�I��H��I��H�)������H��ЃE��}�~��E��}��o�����H��0[A_]���UH��AWSH��@��H�����I�[�      Lۉ}̉uȉUĉM�L�E��E���� �E�``` �E���� �EĉE��ẺE܋E��E؋EȉEԋE؍P��E��xH�M��E�I��A�    �   ��I��H�J������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H�J������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H�J������H��ЋEԍP��E܍pH�M��E�I��A�    �Ѻ   ��I��H�J������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H�J������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H�J������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H�J������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H�J������H��ЋEԍP��E܍p�M��E�ȃ�H�M�I��A�    �Ѻ   ��I��H�J������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H�J������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H�J������H��ЋE؍P��M܋E�ȍp��E���H�M�I��A�    �   ��I��H�J������H��АH��@[A_]���UH��AWSH����H�����I�)�      Lۉ}�H�u�H�E�� ��H�E��@9�sH�E��P#H�E��@9�r"H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@��u)H���������H�H��E�H�։�H��0������H���H�E�H�PH�E��@#��H�H�E�H�PH�E�H�@�U�H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  H�E��@��u0H���������H�H� H��t�E�����I��H�q#������H��ЋE�H��[A_]���UH��H����H�����I���      L�H�}��E�    H�E�@��u]H�E�@'�PH�E�P'��H�E�P#H�E�@'9�r�H�E�H�PH�E�@'��H��H�H�E�H�PH�E�H�@� ���E��   H�E�@��tH�E�@��uiH�E�@#��u������ZH�E�P'H�E�@#9�r������AH�E�H�PH�E�@'��H�H�E�H�PH�E�H�@� ���E�H�E�@'�PH�E�P'�E�����UH��H����H�����I���      L�H���������H�H� H�E��E�    H�E��@��uWH�E��P#H�E��@'9�w�    �AH�E�H�PH�E��@'��H�H�E�H�PH�E�H�@� ���E�H�E��@'�PH�E��P'�E�����UH��H����H�����I��      L�H���������H�H� H�E��E�    H�E��@��uXH�E��@'�PH�E��P'��H�E��P#H�E��@'9�r�H�E�H�PH�E��@'��H��H�H�E�H�PH�E�H�@� ���E��E�����UH��AWH��(��H�����I�a�      L�H�}�H�u�H�U����u�    �(H�M�H�U�H��H��I��H�hL������H���H�E�H�E�H��(A_]���UH��AWSH�� ��H�����I���      L�H�}�H�}� u
������   H�}� tH�E؋@����tH�E��@"<t������zH�E؋@%�   ��u�    �cH�E؋@#H�U؋J�    ��E�H�E؋@��@��u�U�H�E؉�H��I��H��V������H���H�E�H��I��H��S������H��ЉE�E�H�� [A_]���UH��AWSH����H�����I�	�      L�H�}�H�}� u������0H�E�H��H�5������H���H�E�H��I��H��T������H���H��[A_]���UH��AWSH�� ��H�����I���      Lۉ}�H�u�H�}� u
�������  H�EЋ@��u
�    �  H�EЋ@��tH�EЋ@��tH�EЋ@��u!H�UЋE�H�։�H��0������H����y  H�EЋ@����unH�EЋP#H�EЋ�+  9�wYH�EЋ�+  ��tKH�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��E�U�H�EЉ�H��I��H��U������H����H�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U܈H�E�� ��H�EЋ@��9�r3H�EЋ@����H�EЉPH�E�f�   H�E�H��H�5������H���H�EЋ@#�PH�EЉP#H�EЋP#H�EЋ�+  9�vH�EЋ�+  �PH�EЉ�+  H�EЋ@���H�EЉP�    H�� [A_]���UH��AWH��(��H�����I�|�      L�H�}�H�}� u
������  H�E؋@��u
�    �v  H�E؋@��tH�E؋@��tH�E؋@��u"H�E�H��H�"2������H��ЉE�E��0  H�E؋P#H�E؋�+  9�r
������  H�E؋@����ulH�E؋P#H�E؋�+  9�wWH�E؋�+  ��tIH�E؋@����H�E؉PH�E؋@#H�U؋r�    ���E�U�H�E؉�H��I��H��U������H���H�E؋@#H�U؋J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@� ���E�H�E�� ��H�E؋@��9�rH�E؋@����H�E؉PH�E�f�   H�E؋@#�PH�E؉P#�E�H��(A_]���UH��SH��H��H�����I���      L�H�}ȉuĉU�H�M�H�}� u�    �y�E�    H�E�H�E��E�    �FH�E�H��H�v8������H��ЉE؃}��u�E�    �u��4H�E�H�PH�U��U؈�E��E��E��E��E�9�w��E�    �u�H��H[]���UH��SH��H��H�����I���      L�H�}ȉuĉU�H�M�H�}� u�    �l�E�    H�E�H�E��E�    �9H�E�H�PH�U�� ���E�H�U��E�H�։�H�Z6������H��ЃE��E��E��E��E�9�w��E�    �u�H��H[]���UH��H����H�����I�:�      L�H�}�H�u��U�}�tZ�}�|�}� t�}�t�nH�E���H�E��P#H�E���H�E��P'�RH�E��@#H�U��H�E��P#H�E��@'H�U��H�E��P'�(H�E���+  H�U�)Љ�H�E��P#H�E��P#H�E��P'�H�E��@#H�U��J�    ��Љ�H�E�f��    ����UH��H����H�����I�\�      L�H�}�H�}� u�    �	H�E��@#������UH��H����H�����I��      L�H�}�H�}� t7H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@����H�E��P������UH��H��(��H�����I���      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H��(��H�����I�]�      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H����H�����I��      L�H�}��E�_   �(�E�Hc�H�E�H�� < u�E�Hc�H�E�H��  �m��}� y����    ����UH��H����H�����I���      L�H�}�H�E�H�E�H�E�H�E��H�E�� </uH�E�H��H�E�H�E�H�E�� ��u�H�E�����UH��H��0  ��H�����I�5�      L�H������H������H������H�E�H������H�E�H������H�E��E�    �?H�E�� ��u�E�Hc�H�E�H��  �H�E�H�PH�U��U�Hc�H�U�H�� ��E��}�_~��E�    �-H�E�H�PH�U��H�E�H�PH�U�� 8�t�   ��E��}�_~͸    ����UH��SH�� ��H�����I�P�      L�H�}�H�u�H�E؋PH�E؋@ЉE�E�H�U����H�8     H�H�¾   H�B=������H��ЉE�}� t
�������   �E�    ��   �E�%�  ��H�8     ��H؋���uf�E�%�  ��H�8     ��H��������E�H�U����H�8     H�H�¾   H��=������H��ЉE�}� t������r�E��m�E�%�  =�  uE�E��E�H�U����H�8     H�H�¾   H�B=������H��ЉE�}� t�������E�H�E؋@$9E����������H�� []���UH��H����H�����I�Ǿ      L؉}��u�H�U�H�M�    ����UH��AWSH��0��H�����I���      Lۉ}�H�u�H�U�H�EȋPH�Eȋ@ЉE�H�Eȋ@ �E܉E�ЉE�   �    H�8     H�<I��H�@v������H����E�    �B�U�E�Љ�H�EЋ ��H�8     H��   H��=������H��ЉE��}� u�E�H�EȋP �E�9�w���H��0[A_]���UH��H����H�����I���      L�H�}�H�u�H�U��R��H�U����H�U�H��H��   I�B=������J� ������UH��AWSH��`��H�����I�D�      L�H�}�H�u�H�U�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�E�H�E�H�E�H��I��H��s������H��ЉE�H�E��@,�E��9  H�E�H�E��H�E�� </uH�E��  H�E��H�E�H�E�� ��u׋U�H�E��@ H�M��	��H�M���H�B=������H��ЉE؃}� t#H�E�H��I��H�[�������H��и    ��   �E�    �f�E���Hc�H�E�H�H�E�H�E��@a��t5H�E��@b����@��t#H�E�H�U�H��H��H��>������H��ЉE���E������}� t�E��}�?~����}� u+�}�?%H�EЋ@k�E�H�E��@ �E؉E�ЉE�m��	�E�    �
�}� �����H�E�H��I��H�[�������H��ЋE�H��`[A_]���UH��AWSH��P��H�����I�/�      L�H�}�H�u�H�U��M�L�E�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�Eغ    �    H��I��H�@v������H��ЋU�H�E��@ H�M��	��H�M؉�H�B=������H��ЉE�}� t#H�E�H��I��H�[�������H��и������   �E�    �T�E���Hc�H�E�H�H�E�H�E��@a��t#H�E�H�U�H��H��H��>������H��ЉE���E������}� t�E��}�?~����}� u:�}�?4�E���Hc�H�E�H�H�EȺ�   H��H��I��H��u������H�����E�����H�E�H��I��H�[�������H��ЋE�H��P[A_]���UH��AWSH��P��H�����I�e�      L�H�}�H�u�H�U�H�E���C  ��u
������	  H�E���C  ��@v/H���������H�<I�߸    H�
�������H��Ҹ������  H�E��PH�E��@ЉE�H�E���?  H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�Eغ    �    H��I��H�@v������H��ЋU�H�E��@ H�M��	��H�M؉�H�B=������H��ЉEԃ}� t!H�E�H��I��H�[�������H��ЋE��  H�E���C  ��H��H��H�E�H�H�E�H�EȺ`   �    H��I��H�@v������H���H�E�H��+H��H�U>������H���H��H�E�H��H��I��H��x������H����E�    �"H�UȋE�H����uH�UȋE�H�� �E��}�_~�H�E��@` H�E���+  H�EȉPo�U�H�E��@ H�M��	��H�M؉�H��=������H��ЉE�H�E�H��I��H�[�������H��ЋE�H��P[A_]���UH��AWSH��`��H�����I��      L�H�}�H�u�H�U��S  I��H���������H���H�E�H�EкS  �    H��I��H�@v������H���H�E��PH�E��@ ��H�EЉP�    I��H���������H���H�U�H�BH�E��PoH�EЉ�+  H�E��PH�EЉ�/  H�E��P H�EЉ�3  H�E��H�EЉ�G  �    I��H���������H���H�U�H��K  H�E�H��K  �    �    H��I��H�@v������H���H�E��@k�E�    I��H���������H���H�E��E������E�    �E�    ��  �   I��H���������H���H�U�H��K  �M�Hc�H��H�H�H�E�H��K  �U�Hc�H��H�H� H�E�H�E��   �    H��I��H�@v������H����E�    �<  H�E��@ �E��H�E��@�H�E��P�E�H�H�4�    H�E�H�ʉH�EЋ�;  �PH�EЉ�;  �E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E�;E�ts�E�H�U����H�U�H��H�¾   H�B=������H��ЉE��}� t:H�E�H��I��H�[�������H���H�E�H��H��T������H��и    �   �E��E�H�E��@�����E�    ��U�E�H��    H�E�HЋ �E�}��u	�E�������E��}��  ������}��t�E��}��  � �����H�E�H��I��H�[�������H���H�E�H��`[A_]���UH��AWSH��p  ��H�����I���      L�H������H�������   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H������H�E�H��H��I��H��q������H���H�U�H�E�H��H��I��H�Kt������H��п�   I��H���������H���H�     H�H�     H���   �    H��I��H�@v������H��п   I��H���������H���H�E�H�EȺ   �    H��I��H�@v������H���H�E�H�E�H�E��   �    H��I��H�@v������H����E�    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ ���    Hǅ���    Hǅ���    Hǅ���    Hǅ ���    Hǅ(���    Hǅ0���    Hǅ8���    Hǅ@���    HǅH���    HǅP���    HǅX���    Hǅ`���    Hǅh���    Hǅp���    Hǅx���    H�E�    H�E�    H������H������H��H��I��H��x������H���������<wt������<au�E�   H�E��@   H�E��     H�U�H�E�H��H��H�OB������H��ЉE�}� t_H�     H�H��I��H�[�������H���H�E�H��I��H�[�������H���H�E�H��I��H�[�������H��и    �  H�E�H�U�H�M�H�E�H��H��H��B������H��ЉE��}� u_H�     H�H��I��H�[�������H���H�E�H��I��H�[�������H���H�E�H��I��H�[�������H��и    �  H�EȋU��P,H�     H�H�M�H�U�H�u�I�ȹ    H��H��D������H��ЉE�}����   �}� tqH�     H�H������H�U�H�u�A�    H��H�}[������H���H�     H�H������H�U�H�u�I�ȹ    H��H��D������H��ЉE�}� ��   H�     H�H��I��H�[�������H���H�E�H��I��H�[�������H���H�E�H��I��H�[�������H��и    ��  �}� t_H�E�H��I��H�[�������H���H�     H�H��I��H�[�������H���H�E�H��I��H�[�������H��и    �r  H�     H�H�U�H�M�H��H��H��H������H���H�E�H�}� ��   H�     H�H��H�E�H��+�`   H��H��I��H��u������H���H�E�H��+H��H��=������H���������<wt������<+t������<au
H�E��@"�H�E��@"H�E��@   H�EȋP,H�E���?  H�     H��PsH�E���C  ������<auH�     H��PoH�E��P#H�E�H��I��H�[�������H���H�     H�H��I��H�[�������H���H�E�H��I��H�[�������H���H�E�H��p  [A_]���UH��AWSH��@��H�����I�E�      L�H�}��   I��H���������H���H�E�H�E�   �    H��I��H�@v������H���H�E�H�E�H�E�   �    H��I��H�@v������H���H�E��@   H�E��     H�U�H�E�H��H��H�OB������H��ЉE܃}� t H�E�H��I��H�[�������H��и�����AH�U�H�M�H�E�H��H��H��F������H��ЉE�H�E�H��I��H�[�������H��ЋE�H��@[A_]���UH��AWSH�� ��H�����I��      L�H�}�H�E�H�@H��I��H�[�������H����E�    �TH�E�H��K  �U�Hc�H��H�H� H��t?H�E�H��K  �U�Hc�H��H�H� H��I��H�[�������H��ЃE��}��  ~���H�E�H��K  H��I��H�[�������H���H�E�H��I��H�[�������H���H�E�    �    H�� [A_]���UH��H�� ��L�����I��      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H�B=������I� ������UH��H�� ��L�����I�:�      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H��=������I� ������UH��AWSH��   ��H�����I�`�      L�H��x���H��p�����l����   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H��x���H�E�H��H��I��H��q������H���H�U�H�E�H��H��I��H�Kt������H��п   I��H���������H���H�E�H�EȺ   �    H��I��H�@v������H���H�E�H�E�H�E��   �    H��I��H�@v������H���H�E��@   H�E��     H�U�H�E�H��H��H�OB������H��ЉE��}� t_H�     H�H��I��H�[�������H���H�E�H��I��H�[�������H���H�E�H��I��H�[�������H��и�����-  H�E�H�U�H�M�H�E�H��H��H��B������H��ЉE��}� u_H�     H�H��I��H�[�������H���H�E�H��I��H�[�������H���H�E�H��I��H�[�������H��и�����  H�EȋU��P,H�EȋPH�Eȋ@ЉE�H�EȋP,H�Eȋ@ �ЋE�ЉE��    I��H���������H���H�E�H�E��    �    H��I��H�@v������H��ЋU�H�Eȋ@ H�M��	��H�M���H�B=������H��ЉE��E�    �E�    �   �E���Hc�H�E�H�H�E��E�;�l���}~H�E��@a��ta�E���Hc�H��p���H�H�E���   H��H��I��H��u������H��ЋE���Hc�H��p���H�H��H��=������H��ЃE����E��}�?�e�����H�E�H��I��H�[�������H���H�E�H��I��H�[�������H���H�E�H��I��H�[�������H��ЋE�H�Đ   [A_]���UH��AWSH��`��H�����I�t�      L�H�}�H�u�H�U�H�M�D�E�H�E�H�E�H�Eغ�   �    H��I��H�@v������H���H�E�H��H�U>������H���H��H�E�H��H��I��H��x������H����E�    �"H�U؋E�H����uH�U؋E�H�� �E��}�_~�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉEп    I��H���������H���H�E�H�EȺ    �    H��I��H�@v������H��ЋU�H�E��@ H�M��	��H�Mȉ�H�B=������H��ЉEă}� t!H�E�H��I��H�[�������H��ЋE���  �E�    �$�E���Hc�H�E�H�H�E�H�E��@a��t�E��}�?~���H�E��@a���G  �}�?�=  �U�H�E؉PsH�E��@a��E���H�E؈PbH�U�H�E�H��H��H��?������H���H�U؉BkH�E؋@k���uOH�E�H��H���������H�<I�߸    H�
�������H���H�E�H��I��H�[�������H��и   ��   �E���@��t$H�E؋@kH�U�H�M�H�Ή�H�fA������H���H�M�H�E຀   H��H��I��H��u������H��ЋU�H�E��@ H�M��	��H�Mȉ�H��=������H��ЉEĐH�E�H��I��H�[�������H��и    �JH�E�H��I��H�[�������H���H�E�H��H��������H�<I�߸    H�
�������H��Ҹ����H��`[A_]���UH��AWSH��P��H�����I��      Lۉ}�H�u�H�U��    I��H���������H���H�E��E�    �E��E��E������E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E��E܋E�;E���   �}� tV�E�H�U����H�U�H��H�¾   H��=������H��ЉẼ}� t#H�E�H��I��H�[�������H��и�����?  �E�H�U����H�U�H��H�¾   H�B=������H��ЉẼ}� t#H�E�H��I��H�[�������H��и������   �E��E�E��E��E�   H�E��@�����E�    ��U�E�EȋE�H��    H�E�HЋ �E�E�H��    H�E�H��     �}��uL�E�H�U����H�U�H��H�¾   H��=������H��ЉE̐H�E�H��I��H�[�������H��ЋE��6�E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��Y���H��P[A_]���UH��AWSH��   ��H�����I���      L�H��h����   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H��h���H�E�H��H��I��H��q������H���H�U�H�E�H��H��I��H�Kt������H��п   I��H���������H���H�E�H�E��   �    H��I��H�@v������H���H��p���H�E�H�E��   �    H��I��H�@v������H���H�E��@   H�E��     H�U�H�E�H��H��H�OB������H��ЉE�}� t<H�E�H��I��H�[�������H���H�E�H��I��H�[�������H��и    ��  H�E�H�U�H�M�H�E�H��H��H��B������H��ЉE��}� u<H�E�H��I��H�[�������H���H�E�H��I��H�[�������H��и�����d  H�E��U��P,H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE��    I��H���������H���H�E�H�E��    �    H��I��H�@v������H��ЋU�H�E��@ H�M��	��H�M���H�B=������H��ЉE�}� tSH�E�H��I��H�[�������H���H�E�H��I��H�[�������H���H�E�H��I��H�[�������H��ЋE��l  �E�    �   �E������E���Hc�H�E�H�H�E�H�E��@a��t!H�E�H�U�H��H��H��>������H��ЉE�}� u9H�E��@a �U�H�E��@ H�M��	��H�M���H��=������H��ЉE�}� ��E��}�?�k����}� tPH�E�H��I��H�[�������H���H�E�H��I��H�[�������H���H�E�H��I��H�[�������H��ЋE��uH�E��@kH�U�H�M�H�Ή�H��^������H��ЉE�H�E�H��I��H�[�������H���H�E�H��I��H�[�������H���H�E�H��I��H�[�������H��ЋE�H�Đ   [A_]���UH��H����H�5����I�a�      Lމ}�E�E��}� u�E��   �E����rH�H     H�H�H     H�����UH��H����H�����I� �      L�H�}��   H�E�H���r�����UH��AWH����H�����I�ř      L�H�8     H�H�U�H�@     H�    H��      �    H�M�   �    H��I��H�@v������H��ѐH��A_]���UH��AWSH��P��H�����I�=�      Lۉ}��u��}� u
�    ��  H�@     H�H=�   v%H�h�������H�<I�߸    H�
�������H��ҐH��      ���u�H��      ��PH��      ��E����E�E�%�  ��t�E��E�    �E�    �E�    �}� t�E��   �E�   �K  �}��  �=  H�8     H�H�E�H�E�    �E�    �  H�E؋@����   H�E؋@9E���   H�E�H�H�E؋@��H�H�E�H�E؋@+E���H�E؉PH�E؋P�E��H�E؉PH�E�H�E�H�8     H�H�E��E�    �mH�E؋@��tH�E��E��WH�E�H�E�H�E�H�E�H�E�H�@H�PH�E�H�PH�E��@   H�E�H�U�H�H�E��U��PH�E�H�U�H�P�E���!�}��   ~��H�E��E��}��   ������E�   ���}� ��   H�8     H�H�E��E�    �~H�E؋@��tH�E��E��hH�E�H�E��E��H��e������H���H�E�H�E�H�U�H��E��E���H�E��PH�E��U��P�E���+E���H�E��PH�E�H�@   ��}��   �u���H��      �    H�@     H�H�PH�@     H�H�E�H��P[A_]���UH��SH��(��H�����I��      L�H�}�H�}� ��  �H��      ���u�H��      ��PH��      �H�E�H�E�H�8     H�H�E��E�    �M  H�E�H� H9E�tH�E��E��2  H�E�H�E�H�@     H�H�P�H�@     H�H�E؋@��uH�E�H��H��e������H����   H�E؋@��uH�E�H�@H�E�H�E�H�@H�P�H�E�H�PH�E�H�@H��tH�E؋@����   H�E�H�@H��uRH�E�H� H��H��e������H���H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    ��}��   �������H��      �    ��H��([]���UH��AWH��H��L�����I��      M�H�}��u�H�E�    �E�    H�}� u�E��   ��H��f������I� ���8  �H��      A� ��u�H��      A� �PH��      A� H�8     I� H�E�H�E�H�E��E�    �   H�E�H� H9E�t
H�E��   H�E�H�E��E�   H�E��P�E��=   v@H�@     I� �U�H�E�H��H���������I�< M�Ǹ    I�
�������M�A����H�E�H� H�E�H�E��P�E��H�E��P�E��}��   �X���H��      A�     �}� u�E��   ��H��f������I� ���H�E�H��HA_]���UH��H�� ��H�����I�v�      L�H�}�H�u��E�    H�E�H�E��   H�E�� ��H�E��@9�sH�E��P#H�E��@9�rH�E��@#    H�E�f�   H�E�H�PH�E��@#��H�H�E�H�PH�E�H�PH�U�H�U�H�R� �H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  �E��}��E����E�����UH��H�� ��H�����I�v�      L�H�}�H�u��E�    H�E�H�E�H�E��@'�PH�E��P'H�E��P'H�E��@9�rH�E��@'   �H�E��P#H�E��@'9�r�H�E��@'�P�H�E��P'�JH�E�H�PH�E��@'��H�H�E�H�PH�E�H�PH�E�H�HH�M���H�E��@'�PH�E��P'�E��}�~��E�����UH��AWSH��0��H�����I���      L�H�}�H���������H�H� H�E�H�E�H�E�H�E�H��I��H��{������H��ЉE�H�E�H��I��H��{������H��ЉE؋U܋E��=   ~
������   H�E�� </uH�E��E�H�HE�H�m�H�E�� </tH�E�H�E�H�PH�U�� /�H�E�H�U�H�E�H��H��I��H��x������H���H�E�H��I��H��{������H��Љ�HE�H�m�H�E�� </u	H�E��  �H�E�H�E��  �    H��0[A_]���UH��AWSH����H�����I�@�      L�H���������H�H� H��I��H��{������H��Ѓ�w
�    �   H���������H�H� H�E�H�E�H��I��H��{������H��Љ�HE��H�E�H�P�H�U��  H�E�� </u�H���������H�H� H��I��H��{������H��Ѓ�vH�E��  �    H��[A_]���UH��AWSH��0��H�����I�T�      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
�    ��  H�E�H��I��H��{������H��ЉE�E�H�H�P�H�E�H�� </u�E�H�H�P�H�E�H��  �}� 
�    �  �}���   H�E�H��� <:u%H�U�H�E�H��H��I��H��x������H����K  H���������H�<I��H�5�������H���H��H�E�H��H��I��H��x������H���H�E�H��I��H��{������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H��x������H����   H���������H�<I��H�5�������H���H��H�E�H��H��I��H��x������H���H�E�H��I��H��{������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H��x������H���H�E�H��0[A_]���UH��H����H�����I��      L�H�}�H�E�H�E�H�}� u�    �+�E�    �H�E�� </u�E�H�E�H�E�� ��u�E�����UH��AWSH��0��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
������   H�E�H��I��H��{������H��ЉE�E�H�HE�H�m��H�E�� </tH�m�H�E�� ��t�E�P��U�����H�E�H�U�H�E�H��H��I��H��x������H���H�E��  �    H��0[A_]���UH��H��8��H�����I���      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �CH�E�H�PH�U�� ���E�H�E�H�PH�U�� ���E�E�+E�E�}� u�}� t
�m��}� u��E�����UH��H��8��H�����I�+�      L�H�}�H�uЉŰẺE�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M����E��P��U���u�H�E�����UH��H�� ��H�����I���      L�H�}���U��E�E��E�H�E�H�E��H�E�H�PH�U��U��m��}� u�H�E�����UH��AWSH��0��H�����I�O�      L�H�}�H�u�H�E�H�E�H�E�H�E��E�    H�E�H�PH�U�� ����I��H��������H��ЉE�H�E�H�PH�U�� ����I��H��������H��ЉEԋE�+EԉE܃}� u�}� t뗋E�H��0[A_]���UH��AWSH����H�����I���      L�H�}�H�u�H�E�H��I��H��{������H��Љ�H�E�H�H�E�H��H��I��H��x������H���H�E�H��[A_]���UH��H�� ��H�����I��      L�H�}�u�H�E�H�E��H�E�� ��9E�uH�E��H�E�H�E�� ��u۸    ����UH��H�� ��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E��3H�E��H�E�� 8�u!H�E�� ��H�E�� ��Ѕ�u�    �'H�E�H�PH�U��H�E�H�PH�U�� 8�t����������UH��H��0��H�����I�"�      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E��  H�E�����UH��AWH��(��H�����I���      L�H�}؉uԋU��҉Uԃ}� uOH�U�H��I��H��{������H��҉�H�E�H���   H�E�� ��tH�E�� ��9E�u	H�E��   H�E�H�E؃�H��űE�i��E�H�E�H�E��H�E�H�E� ������H�E� ��!�%������u%H�E� 3E䍐����H�E� 3E���!�%������t�H�E�H�E��H�E�H�E�� ��tH�E�� ��9E�u�H�E�H��(A_]���UH��H��@��H�����I�|�      L�H�}�H�u�H�U�H�U�H�U������   H�U�H�������   H�E�    H�E�    H�E�    H�E�    �H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�t�H�E�H+E��'H�U����H�Uȉ�H��H�My������H���H+E�����UH��H����H�����I�F�      L�H�}�H�E�H�E��H�E�H�E�� ��u�H�E�H+E�����UH��AWSH��@��H�����I���      L�H�}�H�u��U�H�E�H�E�H�E�H�E��E�    �kH�E�H�PH�U�� ����I��H��������H��ЉE�H�E�H�PH�U�� ����I��H��������H��ЉEԋE�+EԉE܃}� u�}� t
�m��}� u��E�H��@[A_]���UH��H��(��H�����I�2�      L�H�}�H�u��U�H�E�H�E�H�E�H�E��}� u)������2H�E�H�PH�U��H�E�H�PH�U�� 8�u�m��}� u����E�����UH��H��8��H�����I���      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �!H�U�H�BH�E�H�E�H�HH�M����E��E�9E�w�H�E��  �E�����UH��AWH����H�����I�3�      L�H�}�H�u�H�M�H�U�H��H��I��H�xz������H��҉�HE�H�E�� ��tH�E���    H��A_]���UH��AWH��(��H�����I���      L�H�}؉u�H�U�H��I��H��{������H��҉E��U�H�E�H�H�E��E�    �H�E�� ��9E�uH�E��H�m��E��E�9E�wڸ    H��(A_]���UH��H��0��H�����I�0�      L�H�}�H�u�H�E�H� H�E�H�}� u�    �vH�E�H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u,�}� u
H�E�    �H�E�H���  H�E�H�U�H�H�E���}� u������UH��H��@��H�����I�s�      L�H�}�H�u�H�E�H�E�H�E�    H�E�    H�E�    H�E�    H�E�� ��u
�    ��   H�E�H��� ��u+�H�E�H�E��H�E�� 8�t�H�E�H+E��   H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�u�H�E�H+E�����UH��H��8��H�����I�@      L�H�}�H�u�H�U�H�}� uH�E�H� H�E�H�}� u
�    ��   �H�E�H�PH�U�� ���E�H�E�H�E��
�E�;E�u��H�E�H�PH�U�� ���E��}� uۃ}� uH�E�H�     �    �   H�E�H��H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u4�}� u
H�E�    �H�E�H��H�E�H�E��  H�E�H�U�H�H�E���}� u������UH��H����H�����I�	~      L�H�}�H�u�H�u�H�M�H��      H�H��H���������H�������UH��AWSH�� ��H�����I��}      L�H�}�H�u�H�E�H��I��H��{������H��ЉE��2�U�H�M�H�E�H��H��I��H�3u������H��Ѕ�uH�E��H�E�H�E�� ��uø    H�� [A_]���UH��AWSH�� ��H�����I�}      L�H�}�H�E�H��I��H��{������H��Ѓ��E�E��I��H���������H���H�E�H�}� u�    �$�U�H�M�H�E�H��H��I��H��u������H��АH�� [A_]���UH��H��8��H�����I�z|      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��U�H�E�H�H�E�H�E�H;E�v[H�E�H;E�sQH�E�H�E��E�HE��H�m�H�m�H�E��H�E��H�E�H;E�u��'H�U�H�BH�E�H�E�H�HH�M���H�E�H;E�u�H�E�����UH��AWH����H�����I��{      L�H�}�H�u�H�M�H�U�H��H��I��H�8x������H���H��A_]���UH��AWH����H�����I�`{      Lډ}�H���������H�<I�׸    H�
�������H�������UH��H����H�����I�{      L؉}��U���H���������H�Hc��������t�E� �E�����UH��H����H�����I��z      L؉}��U���H���������H�Hc��������t�m� �E�����UH��AWSH��0��H�����I�ez      L�H�}ȉuĉU��M��U�H�E�H��H���������H�<I�߸    I�
�������I�A��H�E�H��I��H���������H���H�E�H�E� �E�H�E� 9E�u��H��0[A_]���UH��AWSH�� ��H�����I��y      L�H�}�H�u�H�E�� ��u�    �LH�E�� <wuH�E�H��I��H���������H���H�U�H�E�H��H��I��H��4������H���H�E�H�E�H�� [A_]���UH��AWH����H�����I�.y      L�H�}�H�U�H��I��H��5������H���H��A_]���UH��AWH����H�����I��x      L�H�}�H�U�H��I��H�5������H���H��A_]���UH��AWH����H�����I��x      L؉}�H�u�H�M��U�H�Ή�I��H�Z6������H���H��A_]���UH��AWSH�� ��H�����I�Dx      L�H�}�H�}� u������VH�E�H��I��H�v8������H��ЉE�H�E؋@��u+H���������H�H��E�H�։�I��H�Z6������H��ЋE�H�� [A_]���UH��AWH����H�����I��w      L؉}�H�u�H�M��U�H�Ή�I��H�Z�������H���H��A_]���UH��AWH����H�����I�Zw      L�H�}�H�U�H��I��H���������H���H��A_]���UH��AWSH��@��H�����I�w      L�H�}ȉu�H�U�H�}� u	H�E��  H�E�H�E�H�E�H�E��E�    H�E�H��I��H�v8������H��ЉEԃ}����   H�E��@��u7�}�u�}� ~+H���������H�H��E�H�։�I��H�Z6������H��Ѓ}�
tk�E�;E�}E�}�u�}� ~H�E�H;E�vH�m��m��:�}��^���H�E�H�PH�U�UԈ�E��D����}�u�}� ~�m���E��)�������}�~	H�E��  ��Eԉ�H�E�H�E�H��@[A_]���UH��AWSH�� ��H�����I��u      L�H�}�H�u�H�}� u�    �^�E�    �2�E�Hc�H�E�H�� ��H�U�H�։�I��H�Z�������H��ЃE�H�E�H��I��H��{������H��ЋU�9�w��E�H�� [A_]���UH��AWH��(��H�����I�u      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I�E:������I�A��H��(A_]���UH��AWH��(��H�����I��t      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I�;������I�A��H��(A_]���UH��AWH����H�����I�Vt      L�H�}�H�U�H��I��H�.a������H���H��A_]���UH��AWH����H�����I�t      L�H�}�H�U�H��I��H��<������H��ҐH��A_]���UH��AWH��(��H�����I��s      L�H�}�H�u��U܋U�H�u�H�M�H��I��H��;������H���H��(A_]���UH��H����H�����I�hs      L�H�}�H�}� u������!H�E��P#H�E���+  9�r�������    ����UH��AWH����H�����I�s      L�H�}�H�U�H��I��H��<������H���H��A_]���UH��AWSH��`  ��H�����I��r      L�H������H������H�������E�    �E�    �  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H���������H���	E�}���  �E�H��    H��h  H�H��h  H�>��H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E��E�H������H�։�I��H�E�������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�}� t(H������H�E�H��H��I��H�>�������H����O  H������H��H��������H�<I��H�>�������H����   H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E�H�������E�H�։�I��H��������H���H������H������H��H��I��H�>�������H����w  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������
   H��H��I��H�}�������H���H������H������H��H��I��H�>�������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������   H��H��I��H�J�������H���H������H������H��H��I��H�>�������H����  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�EȾ   H��fHn�I��H�8�������H���H������H������H��H��I��H�>�������H����]  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eк
   H��H��I��H���������H���H������H������H��H��I��H�>�������H����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ
   H��H��I��H�}�������H���H������H������H��H��I��H�>�������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ   H��H��I��H�}�������H���H������H������H��H��I��H�>�������H����G  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�E�   H��fHn�I��H�8�������H���H������H������H��H��I��H�>�������H����   H������H�ƿ%   I��H�E�������H��ЋE�Hc�H������H�� ��H������H�։�I��H�E�������H����4�E�Hc�H������H�� ��H������H�։�I��H�E�������H��ЃE��E�Hc�H������H�� ��������    H��`  [A_]���UH��H����H�����I�3j      L؉��E��E�    �E��S��%wa��H��    H��a  H�H��a  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��i      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H�0�������L��Љ�<�����<���H���   A_]���UH��H�� ��H�����I��h      L�H�}�H�u�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E�����UH��AWSH��  ��H�����I�,h      L�H������H������H��x����E�    H������H�E�f�E�  �E� �E�    �/  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H���������H���	E܃}���  �E�H��    H�R`  H�H�G`  H�>��H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E��E�H�U�H�E�H��H��H�V�������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H�}� t'H�U�H�E�H��H��H�V�������H���H�E��e  H�E�H��������H�4H��H�V�������H���H�E��7  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E�H�������E�H�։�I��H��������H���H������H�E�H��H��H�V�������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������
   H��H��I��H�}�������H���H������H�E�H��H��H�V�������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������   H��H��I��H�J�������H���H������H�E�H��H��H�V�������H���H�E��3  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�E��   H��fHn�I��H�8�������H���H������H�E�H��H��H�V�������H���H�E��x  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�E��
   H��H��I��H���������H���H������H�E�H��H��H�V�������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ
   H��H��I��H�}�������H���H������H�E�H��H��H�V�������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ   H��H��I��H�}�������H���H������H�E�H��H��H�V�������H���H�E��e  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�Eо   H��fHn�I��H�8�������H���H������H�E�H��H��H�V�������H���H�E��   H�E�H��������H�4H��H�V�������H���H�E�fǅ����  �E�Hc�H������H�� ������H������H�E�H��H��H�V�������H���H�E��8�E�Hc�H������H�� �E�H�U�H�E�H��H��H�V�������H���H�E��E��E�Hc�H������H�� �������H�E��  H�U�H������H)�H��H�Ā  [A_]���UH��H����H�����I�]_      L؉��E��E�    �E��S��%wa��H��    H��X  H�H��X  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��^      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H�������L��Љ�<�����<���Hc�H�����H��  ��<���H���   A_]���UH��AWH���   ��L�����I��]      M�H����������H�����H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H����������H�����H��M��H�/�������L��Љ�<�����<���H���   A_]���UH��AWSH��0��H�����I��\      L�H�}؉u�H�U�H�M��}�   v
�    �   H�U�H�E�H��H��      H�<I��H�������H��ЉE�}���  ~�   �I�E�E�}� ~:�U�H�E�H��      H�4H��I��H��u������H��ЋE�Hc�H�E�H��  �E�H��0[A_]���UH��AWH����H�����I��[      L؉}�H���������H�H�
�U�H�Ή�I��H�Z�������H���H��A_]���UH��AWSH�� ��H�����I��[      L�H�}�H�}� tj�E�    �?H���������H�H��E�Hc�H�E�H�� ��H�։�I��H�Z�������H��ЃE�H�E�H��I��H��{������H��ЋU�9�w���H�� [A_]���UH��AWH���   ��L�����I��Z      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H�0�������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I��Y      M�H��8���H��0���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�H��������I�<M�׸    H�
�������L�������UH��AWH����H�����I�RY      L�H�}�H�U�H��I��H�d�������H��ҐH��A_]���UH��AWH��(��H�����I�Y      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H��������H��Ѹ    H��(A_]���UH��AWH��(��H�����I��X      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H��������H����H�E�H�E�� < tH�E�H   H9E�sH�E�� <
u�H�E��  H�E�H;E�����H��(A_]���UH��AWSH��0��H�����I��W      L�H�}�H�uЉỦM�H��     H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H��������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H��     H�H�E�H��     �0H��     �D �}�u-�U�H�E�    H��I��H���������H���H�U�H��   �}�u+�U�H�E�    H��I��H�ֺ������H��Љ�H�EЉ�[�}�u,�U�H�E�    H��I��H�ֺ������H��Љ�H�E�f��)�U�H�E�    H��I��H�ֺ������H��Љ�H�EЈ�    H��0[A_]���UH��AWSH��0��H�����I�ZV      L�H�}�H�uЉỦM�H��     H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H��������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H��     H�H�E�H��     �0H��     �D �}�u'H�E�H��I��H�#�������H����Z�H�E�� �+�}�u%H�E�H��I��H�#�������H���fH~�H�U�H��    H��0[A_]���UH��SH��8��H�����I�U      L�H�}�H�u�H�U��E�    �E�    ��  �E�    �E�Hc�H�E�H�� ������%��  �E��E�Hc�H�E�H�� ������lu�E��E�   �E�Hc�H�E�H�� ����H�0�������H���	E�}��o  �E�H��    H�tO  H�H�iO  H�>��H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H��������H�����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H�Q�������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H����?  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��������H�����   H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��������H����jH�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H������E��E�Hc�H�E�H�� ��������E�H��8[]���UH��H����H�����I��P      L؉��E��E�    �E��S��%wa��H��    H�cL  H�H�XL  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I�P      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H�Ԫ������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I�*O      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H�Ԫ������L��Љ�<�����<���H���   A_]���UH��H����H�����I�:N      L؉}�H�u�H�}� u������w�}��u������jH�E��@#��tH�E��@#�P�H�E��P#H�E��@#H�U��J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U���E�����UH��AWSH����H�����I��M      L�H���������H�H� H��I��H�v8������H��ЉE�}��t+H���������H�H��E�H�։�I��H�Z6������H��ЋE�H��[A_]���UH��AWH��(��H�����I��L      L�H�}�H�u�H�U�H��������H�<I�ϸ    H�
�������H�������UH��H����H�����I��L      L�H�}��	   H�E�H���r�����UH��SH����H�����I�hL      L�H�}�H�}� u.H��     H�<H�R�������H���H��     H��H�E�H��H�R�������H���H�E�H��[]���UH��AWSH��0��H�����I��K      L�H�}�H�u�H�E�H�"�������H�4H��I��H�.�������H���H�E�H�}� u
������   �E�    H�E�H��I��H��{������H��ЉE܃}�`~	�E�   �$H�E�H�P+H�E�H��H��I��H��x������H���H�E��@���H�E��PH�E�H��I��H�Ć������H��ЋE�H��0[A_]���UH��H��0��H�����I��J      L؉}�H�u�H�E�H�E��E܉E��E�    �}� y,H�E�H�PH�U�� -�}�   �u�E�����E���E��؉E�H�E�H�E�M�Hc�Hi�gfffH�� ��������)�����)��ʉЍH0H�E�H�PH�U�ʈ�E�Hc�Hi�gfffH�� ����)ЉE�}� u��}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWSH��@��H�����I��I      L�H�}�H�u��U�H�}� u#H�E�H�E�H�E�H�PH�U�� 0H�E��  �  H�E�H�E؋E�Hc�H�E�H�H�E��3H�E؃��E�H�m��}�	~�7   ��0   �U��H�m���H�E�H�E�H;E�wËE�Hc�H�E�H��  H�E�H�E��E�    �8H�E�� <0uH�E��"H�U�H�E�H��H��I��H��x������H�����E��E�;E�|�H�E�H�E�H�E�H��I��H��{������H��Љ�H�E؋E�H�U�)Љ�H�M�H�E�HȾ    H��I��H�@v������H���H��@[A_]���UH��AWH����H�����I�3H      L؉}�U�    ��I��H��f������H���H��A_]���UH��AWH����H�����I��G      L؉}�u�U��U��I��H���������H���H��A_]���UH��AWH����H�����I��G      L�H�}�H�U�H��I��H��i������H��ҐH��A_]���UH��AWH����H�����I�KG      L�H�}�u�M�H�U��H��I��H��k������H���H��A_]���UH��H����H�����I��F      L؉}�u�E��}�E��E��}�ЉE��}� x�E���y�E����E��E�+E�E��!�}� y�E���~�E����E��U��E�ЉE�H�E�����UH��H�� ��H�����I�rF      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H�� ��H�����I��E      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H��H��H�����I�E      L�H�}�H�u��U�H�E�H�E�H�E�H�PH�U�� ���E�E���H���������H�H������ ��uǃ}�-u�E�   H�E�H�PH�U�� ���E��"�E�    �}�+uH�E�H�PH�U�� ���E�}� t�}�u9�}�0u3H�E�� <xtH�E�� <XuH�E�H��� ���E�H�E��E�   �}� u�}�0u�   ��
   �E��}� t	H��   ������H�E�E�Hc�H�E�H�H��H�ЉE؋E�Hc�H�E�H�H��H�E�}� t�}� ~�E�)E�H�E��]�H�E�    �E�    �E���H���������H�H��������t�m�0�[�E���H���������H�H���������5  �E���H���������H�H��������t�7   ��W   )E�E�;E���   �}� ��   �}� tgH�E�H;E�|H�E�H;E�u0�E�;E�~(�E�����H�E�   �H���������H�� �����   �E�   �E�H�H�U�H��H�E��E�H�H)E��eH�E�H;E�H�E�H;E�u-�E�;E�~%�E�����H�E����H���������H�� �����$�E�   �E�H�H�U�H��H�E��E�H�HE���H�E�H�PH�U�� ���E��y������H�}� t�}� t
H�E�H���H�E�H�U�H�H�E�����UH��AWH����H�����I��A      L�H�}�H�M�
   �    H��I��H�ֺ������H���H��A_]���UH��AWH����H�����I��A      L�H�}�H�M�
   �    H��I��H�ֺ������H���H��A_]���UH��AWAVAUATSH����H�����I�9A      L�H�}�H�uȉU�L�eп    L��L�`� �؉���H���������H�H������ ��uЃ�-u�   L��L�`� �����+uL��L�`� �؃}� t�}�u-��0u(A�$<xt	A�$<XuI�D$� ��I���E�   �}� u��0u�   ��
   �EċE�Hc������    H��I�ǋE�Hc������    H��H�Љ�A�    A�    ����H���������H�H��������t��0�T����H���������H�H��������tz����H���������H�H��������t�7   ��W   )�;]�}GE��x
M9�wM9�u��9�~A������A�   �E�H�L��Hc�I�L��L�`� ���;������E��yA�����H���������H�� "   �	����tI��H�}� tE��tI�D$��H�E�H�U�H�L��H��[A\A]A^A_]���UH��H����H�����I��>      L؉}��   �   ���r����UH��AWSH����H�����I��>      L�H�}�H�E�H�%�������H�4H��I��H�8x������H��Ѕ�uH���������H�H� ��    H��[A_]���UH��AUATSH�� ��H�����I�C>      L�H�}�H�u�H�`     ��E�L�e�H�]�E�,$L��L�`��H��H�XD�(�m��}� uې�H�� [A\A]]���UH��H��8��H�����I��=      L�H�}�H�u�H�U�H�`     ��E�H�E�H�E�H�E�H�E�H�E�H�E�H�E�� ���E�H�E�H�PH�U�H�U���H�E�H�PH�U�H�U���H�E�H�PH�U��U���m��}� u�������UH��SH��H��H�����I�=      L�H�}�H�u�H�`     ��E�H�E�H+E��EȋE�9E���  �E�����EȺ    ��E��EȋU�H�E�H�H�E�H�E�H�E�H�E�H�E�E�H�H��H��H�E�H�H�E�H�E�H;E�sjH�X     H�H�U�H�E�H��H���щEă}� u/�E�H�H��HE�H�U�H�E�H��H��H���������H�����  �}� y�E�H�HE���  �H�E�H;E���   H�X     H�H�U�H�E�H��H���щEă}� u)�E�H�HE�H�U�H�E�H��H��H���������H���뢃}� ��   H�E�H;E�uA�E�H�HE�H�U�H�M�H�E�H��H��H�'�������H��ЋE�H�HE�H�E�H�E��M���H�U�H�E�H��H��H���������H��ЋE�H�H��HE��E�H�HE���   �E�H�H��HE�����H�E�H;E���   H�E�H+E�H��H�E�H+E�H9�|4�E�Hc�H�E�H�H�E�H��H��H���������H���H�E�H�E������H�U�H�E�H��H��H���������H��ЋE�Hc�H�E�H�H�E������E�H�H��HE�H�U�H�M�H�E�H��H��H�'�������H��ЋE�H�H��HE�H�E�H�E������H��H[]���UH��H�� ��H�����I�-:      L�H�}��u�U�H�M�H�X     H�U�H��U�H�`     ��U��U���H�U�H�H�U�H��H��H���������H��А����UH��AWH����H�����I��9      L�H�}�H�)�������H�<I�׸    H�
�������H��Ѹ����H��A_]���UH��H��@��H�����I�P9      L�H�}�H�u�H�U�H�U��H�E�H�U����H���������H�Hc���҃� ��u��E�    H�U���҃�+t��-u�E�   H�E�H�H���������E��E�    �E�    �E�    �;�M�H�P���������Y�H�U���҃�0�*��X��E�H�E��E�H�U����H���������H�Hc���҃���u�H�U����.uuH�E��?�M�H�P���������Y�H�U���҃�0�*��X��E�H�E��E��E�H�U����H���������H�Hc���҃���u��U�)U�}� uH�H�������f���  �}� t�E�H�X�������f(fW��E�H�U����etH�U����E��   �E�    H�E�H�U���҃�+t��-u�E�   H�E��E�    �%�M܉����҉�H�U���҃�0ʉU�H�E�H�U����H���������H�Hc���҃���u��}� t�U�)U���U�U�}����|	�}�   ~H�����������   H�P���������E��E�E܃}� yF�]��A�E܃���t&�}� y�E��^E��E���E��YE��E��}��E��Y��E��}� u�H�}� tH�E�H�U�H��E�����UH��H����H�����I�6      L؉}�H�E�   �E�    �H�U�H��H��H�H�H�E��E��E�;E�|�H�E�����UH��AWSH��@��H�����I��5      L��E�H�}��u�H�}� u	H�E��  H�E�H�E�H�p�������f��f/E�v,H�E�H�PH�U�� -�E�H�x�������f(fW��E��E�H���������f/s�E��H,�H�E��/�E�H�����������\��H,�H�E�H�       �H1E�H�E�H�E�H�E�H��x�H*��H��H���H	��H*��X��M��\�f(��EȋE���H���������H���H��x�H*��H��H���H	��H*��X��YE�H���������f/s�H,�H�E��*H�����������\��H,�H�E�H�       �H1E�H�E�H�E�H�M�H�U�H�E�H�h�������H�43H��I�߸    I�A�������I�A��H�E�H��@[A_]���UH��AWH����H�����I��3      L�H�}�H�U�    H��I��H���������H���H��A_]���UH��AWH����H�����I�3      L�H�}�H�u�H�M�H�U�H��H��I��H���������H����Z�H��A_]���UH��AWH��(��H�����I�%3      L�H�}�H�u�H�M�H�U�H��H��I��H���������H����E��E�H��(A_]���UH��H����H�����I��2      L؉}��E����3E�)�����UH��H��@��H�����I��2      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�    H�}� y>H�E�H�PH�U�� -H�       �H9E�uH��������H�E�H�E��H�E�H��H�E�H�E�H�E�H�M�H�gfffffffH��H��H��H��H��?H)�H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U��ʈH�M�H�gfffffffH��H��H��H��H��?H)�H��H�E�H�}� u�H�}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U߈H�E�H;E�w�H�E�����UH��AWH��8��H�����I�1      L�H�}�H�uЉU�H�U�H�U�H�}� yH�U�H�JH�M��-H�]�H�U�H�U��}�u$H�M�H�u�   H��I��H�J�������H����H�M�H�U�H��H��H�_�������H���H�E�H��8A_]���UH��H��0��H�����I�p0      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E�H�M�H���������H��H��H��H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U�ʈH�E�H���������H��H��H��H�E�H�}� u�H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWH��8��H�����I�u/      L�H�}�H�uЉU�H�U�H�U�H�U�H�U��}�u$H�u�H�M�   H��I��H�J�������H����H�M�H�U�H��H��H���������H���H�E�H��8A_]���UH��H����H�����I��.      L؉}������UH����H�����I��.      Lظ   ]���UH��H����H�����I��.      L�H�}��    ����UH��H����H�����I�b.      L�H�}�H���������H�H� ����UH��H����H�����I�'.      L�H�}�H���������H�H� ����UH��H�� ��H�����I��-      L�H�}��u�H�U�H�M�    ����UH����H�����I��-      Lظ    ]���UH��H����H�����I��-      L��E�H���������f������UH��H����H�����I�R-      L��E�H���������f������UH��H����H�����I�-      L��E��}�H���������f������UH��H����H�����I��,      L��E�H�}�H���������f������UH��H����H�����I��,      L��E��M�H���������f������UH��H��(��H�����I�b,      L��E��M��E��U��U��E��E��E������������������������������]��E�����UH��H����H�����I��+      L��E����E����]��E�����UH��H����H�����I��+      L��E�H���������f������UH��H����H�����I��+      L��E�H���������f������UH��H����H�����I�G+      L��E�H���������f������UH��H����H�����I�+      L��E�H�����������E��E�����UH��H����H�����I��*      L��E�H���������f������UH��H����H�����I��*      L��E�H���������f������UH��H����H�����I�X*      L��E�H���������f������UH��H����H�����I�*      L��E�H���������f������UH��AWH����H�����I��)      L��E��E�H���������H�f(�fHn�I��H���������H���H��A_]���UH��H����H�����I��)      L؉}�H�u�    ����UH��AWH����H�����I�Q)      Lډ}�H�u�H���������H�<I�׸    H�
�������H�������UH��AWH��(��H�����I��(      Lى}�H�u�H�U�H���������H�<I�ϸ    H�
�������H�������UH��AWSH�� ��H�����I��(      L�H�}�H��������H�<I�߸    H�
�������H����E�    �.�E�H�H��    H�E�HЋ ��I��H��������H��ЃE��}�?~̸����H�� [A_]���UH��AWH����H�����I�
(      L�H�}�u�H��������H�<I�׸    H�
�������H�����f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     @                                                                     ~ � � � � � � � � ~             ~ � � � � � � � � ~                 l � � � � | 8                   8 | � | 8                   < < � � �   <                < ~ � � ~   <                      < <              � � � � � � � � � � � � � � � �           < f B B f <           � � � � � � � � � � � � � � � �        2 x � � � � x             < f f f f <  ~               ? 3 ? 0 0 0 0 p � �              c  c c c c g � � �               � < � < �             � � � � � � � � � � �               > � >                  < ~    ~ <                f f f f f f f   f f              � � � {                | � ` 8 l � � l 8  � |                       � � � �              < ~    ~ <  ~              < ~                           ~ <                      �                         0 ` � ` 0                         � � � �                       ( l � l (                      8 8 | | � �                   � � | | 8 8                                                 < < <                  f f f $                             l l � l l l � l l           | � � � |   � � |               � �   0 ` � �             8 l l 8 v � � � � v           0 0 0 `                             0 0 0 0 0 0               0         0                   f < � < f                         ~                                    0                     �                                                           0 ` � �             8 l � � � � � � l 8              8 x       ~             | �    0 ` � � �             | �   <    � |               < l � �                 � � � � �    � |             8 ` � � � � � � � |             � �     0 0 0 0             | � � � | � � � � |             | � � � ~     x                                                       0                  0 ` 0                      ~     ~                     ` 0      0 `             | � �                       | � � � � � � � |              8 l � � � � � � �             � f f f | f f f f �             < f � � � � � � f <             � l f f f f f f l �             � f b h x h ` b f �             � f b h x h ` ` ` �             < f � � � � � � f :             � � � � � � � � � �             <         <                   � � � x             � f f l x x l f f �             � ` ` ` ` ` ` b f �             � � � � � � � � � �             � � � � � � � � � �             | � � � � � � � � |             � f f f | ` ` ` ` �             | � � � � � � � � |           � f f f | l f f f �             | � � ` 8   � � |             ~ ~ Z       <             � � � � � � � � � |             � � � � � � � l 8              � � � � � � � � � l             � � l | 8 8 | l � �             f f f f <     <             � � �   0 ` � � �             < 0 0 0 0 0 0 0 0 <               � � � p 8                 <         <          8 l �                                                   �       0                                     x  | � � � v             � ` ` x l f f f f |                   | � � � � � |                < l � � � � v                   | � � � � � |              6 2 0 x 0 0 0 0 x                   v � � � � � |  � x       � ` ` l v f f f f �                 8      <                        f f <       � ` ` f l x x l f �             8         <                   � � � � � � �                   � f f f f f f                   | � � � � � |                   � f f f f f | ` ` �             v � � � � � |                � v f ` ` ` �                   | � ` 8  � |              0 0 � 0 0 0 0 6                    � � � � � � v                   � � � � � l 8                   � � � � � � l                   � l 8 8 8 l �                   � � � � � � ~   �             � �  0 ` � �                 p                                        p         p                       v �                        8 l � � � �                               ��� ��� ~~~                                 uuu ��� ��� ���                                 ��� ��� ��� ��� ;;;                          ��� ��� ~~~ ��� ���                         ��� ��� ���     ��� ���                         ��� ���      ��� ��� ppp                 @@@ ��� ���         III ��� ���                 ��� ��� ��� ��� ��� ��� ��� ���                 ��� ���                 zzz ��� ���         ``` ��� ���                     ��� ���         ��� ��� MMM                     ��� ��� bbb     ��� ���                         ||| ��� ���      ��C? This help cd Change current directory clear Clear screen copy Copy file or directory date Date del Delete file or directory dir List directory echo This --- exit Exit shell help info This System information mov Move file or directory new New file or directory reboot Reboot system rename Rename file or directory poweroff Turn off the computer time Time version Shell version PWD <%s> ~ $ %s  %s: command not found
 ./ Function not implemented
 rename: error
 w Sirius OS (Kernel mode: AMD64 or x86_64)
CPU: %s
 Commands:
    Erro, arquivo ou directorio nao encontrado
 .. %s/.     cd: %s: No such file or directory
 ./ dir: error
 dir: empty
 %s
 BitMAP error
 Not suport BitMAP 4-bit Not suport BitMAP > 8-bit       Entrada maior que o limite
 Erro ao criar o arquivo "%s"
       Error ao criar o arquivo "%s", atingio o limite de arquivos na entrada de directorio
   Panic: __malloc, sem espaco na tabela de alocacao
      panic: realoc sem espaco, %lx size = %d %d
 PWD strerrorr
                              (((((�AAAAAABBBBBB                                �Dubug: %s %x %x
        (null)  ����������������������Y����������������������`�������`�������������������������������������������������������������������������������������������Λ��������������2�������2�������P���������������������������������������k���������������������������������������������������������������������������������������G�������Y���������������}�������t���������������Y�������������������������������������������������������������������������������P���������������b�����������������������k�������(null) %        ����������������J����������������������[�������	�������	�����������������������������������������������������������������������������������������������ģ������u�������&�������ץ������ץ������&�������\�������\�������\�������\�������A�������\�������\�������\�������\�������\�������\�������\�������\�������\�������\��������������/�������\�������S�������J�������\�������/�������\�������\�������\�������\�������\�������\�������\�������\�������\�������&�������\�������8�������\�������\�������A�������panic: sscanf()
        ����������������������g�������ӱ�������������?�������?��������������������������������������������������������������������������������������������������������������������������������������������������������������ҳ����������������������������������������������������������������������������������������������������������۳���������������������������������������������������������������������������������������������������ɳ��������������������ҳ������panic: freopen()
 r+ PWD call system funtion error. 
                 $@       �        %lu.%lu                �              �C                                                                        �_�
�@panic: signal()
 panic: sigaction()
 panic: setjmp()  panic: longjmp                                                                                                                                                                                                                                                                                                                                                                                    �$ �     �     �   �. �   �$ �   �. �   �$ �      �   �$ �      �   ` �   % �   (% �                           h �   9,  �   j �   t �   X0  �   w �   � �   �/  �   � �   � �   �/  �   � �   � �   </  �   � �   � �   ~.  �   � �   � �   -.  �   � �   � �   �-  �   � �    �   �-  �    �    �   9,  �   j �    �   �+  �   ! �   9 �   B+  �   = �   T �   �*  �   X �   n �   `*  �   u �   � �   �)  �   � �   � �   �)  �   � �   � �   &)  �   � �   � �   �(  �   � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          zR x�  ,      @����   E�CG����B�A�          L   ����<    E�Cs�  $   l   ����    E�CG��{�B�A�(   �   n����   E�CG��x�B�A�      �   �����    E�C��    �   n���z   E�CG��         ����Z    E�CF�J�A�    $  ����Z    E�CF�J�A�   H  4���@    E�Cw�  $   h  T����    E�CG����B�A�   �  ����@    E�Cw�  $   �  �����    E�CG����B�A�    �  f���Z    E�CF�J�A�$   �  �����    E�CJ����B�A�(   $  ���h   E�CG��U�B�A�      P  M���2    E�Ci�      p  _���Z    E�CF�J�A�    �  ����Q    E�CF�A�A�$   �  �����    E�CG����B�A�    �  X���Z    E�CF�J�A�      ����Z    E�CF�J�A�    (  ����h    E�CF�X�A�,   L  ���'   E�CG���B�A�       ,   |  ����   E�CG����B�A�          �  � ���    E�C�� $   �  W��   E�CE��A�   $   �  D���    E�CG����B�A�$     ����    E�CG����B�A�(   D  j���   E�CG����B�A�   (   p  ���j   E�CG��W�B�A�       �  &���    E�CE���� (   �  ���   E�CG���B�A�       �  ����    E�CE���� (     I���   E�CG��q�B�A�   $   <  ���   E�CG����B�A�   d  ���9    E�Cp�     �  ���+    E�Cb�     �  ����    E�C��     �  ���   E�CE����   �  ���I    E�C@�       ���u    E�CE�f�A�(   ,  -���   E�CG����B�A�   (   X  ����   E�CG����B�A�   $   �  ����    E�CG����B�A�,   �  N��2   E�CG���B�A�       (   �  P��Z   E�CG��G�B�A�        ~��   E�C�   (  |���    E�C��    H  ���    E�C��     h  ���p    E�CF�`�A�$   �  ����    E�CG����B�A�$   �  ���r    E�CG��_�B�A�(   �  ���   E�CG��	�B�A�   $     � ���   E�CF���A�       0  y"���    E�CE���A�    T  #���    E�CE���A�   x  �#���    E�C��    �  d$��A    E�Cx�      �  �$��i    E�C`�        �  �$��U    E�CL�    �  �$��U    E�CL�    	  4%��i    E�C`�    <	  }%��g    E�C^�    \	  �%���    E�C�� $   |	  �&���   E�CE�{�A�      �	  �'��9    E�Cp�  $   �	  (���    E�CG����B�A�   �	  �(��^    E�CU� (   
  )��   E�CG���B�A�   (   8
  �*���   E�CG����B�A�   (   d
  �,��]   E�CG��J�B�A�   (   �
  �.��   E�CG��l�B�A�   (   �
  2��D   E�CJ��.�B�A�   (   �
  (9��:   E�CG��'�B�A�   $     6:��    E�CG����B�A�   <  ;���    E�C��    \  �;���    E�C�� (   |  v<���   E�CJ����B�A�   (   �  9@��i   E�CG��V�B�A�   (   �  vC��H   E�CG��5�B�A�   (      �E��e   E�CJ��O�B�A�      ,  �I��a    E�CX�    L  J��9    E�Cp�      l  %J���    E�CF�w�A�(   �  �J��'   E�CG���B�A�   $   �  �M��   E�CE���A�   $   �  \O���   E�CF���A�        �P��    E�C��    ,  �Q���    E�C�� (   L  zR��O   E�CG��<�B�A�   $   x  �S���    E�CG����B�A�(   �  aT��C   E�CG��0�B�A�      �  xV��k    E�Cb� $   �  �V���    E�CG����B�A�     �W���    E�C��    4  �W��w    E�Cn�    T  PX��b    E�CY� $   t  �X���    E�CG����B�A�$   �  %Y��z    E�CG��g�B�A�   �  wY��a    E�CX�    �  �Y���    E�C��      2Z��{    E�Cr� $   $  �Z��+   E�CF��A�      L  �[��6   E�C-�   l  �\��L    E�CC� $   �  �\���    E�CG����B�A�   �  r]���    E�Cw�    �  �]��}    E�Ct� $   �  /^��r    E�CF�b�A�    $     y^���    E�CF���A�       D  �^���    E�C��    d  �_��3   E�C*�   �  �`��7   E�C.�   �  �a��W    E�CN� $   �  �a���    E�CG����B�A�$   �  Rb���    E�CG����B�A�     �b���    E�C�� $   4  lc��V    E�CF�F�A�       \  �c��P    E�CF�       |  �c��U    E�CL�    �  �c��U    E�CL� $   �  4d���    E�CG����B�A�$   �  �d���    E�CG����B�A�$     e��K    E�CF�{�A�     $   4  ?e��K    E�CF�{�A�     $   \  be��S    E�CF�C�A�    $   �  �e���    E�CG����B�A�$   �  �e��S    E�CF�C�A�    $   �  (f��K    E�CF�{�A�     ,   �  Kf��[   E�CG��H�B�A�       $   ,  vg���    E�CG����B�A�$   T  �g��]    E�CF�M�A�    $   |  'h��]    E�CF�M�A�    $   �  \h��K    E�CF�{�A�     $   �  h��L    E�CF�|�A�     $   �  �h��Y    E�CF�I�A�         �h��Y    E�CP� $   <  i��K    E�CF�{�A�     (   d  0i���   E�CJ��{�B�A�       �  �q���    E�C��     $   �  r���    E�CI���A�       �  �r��l    E�Cc� (   �  *s���   E�CJ����B�A�       (  �{���    E�C��     $   L  Y|��   E�CI���A�    $   t  2}���    E�CI���A�    $   �  �}���    E�CG����B�A�$   �  �~��\    E�CF�L�A�    $   �  �~���    E�CG����B�A�$     Z���    E�CI���A�       <  '����    E�CI�    $   \  ����L    E�CF�|�A�         �  ̀��e    E�CF�U�A�    �  ����    E�CF���A�(   �  �����   E�CG����B�A�   (   �  ���=   E�CG��*�B�A�   $   $  ���\   E�CE�M�A�      L  H����    E�C�� $   l  ҈���    E�CI���A�    $   �  �����    E�CI���A�       �  b����    E�C�� $   �  ����    E�CG��z�B�A�     Y���Y    E�CF�       $  ����9    E�Cp�  $   D  �����    E�CE�q�A�    $   l  ����    E�CG����B�A�   �  ӌ��G   E�C>�,   �  ����u   E�CG��b�B�A�       $   �  ?���M    E�CF�}�A�     $     d���O    E�CF��A�     $   4  ����L    E�CF�|�A�     $   \  ����S    E�CF�C�A�       �  ڏ���    E�C�    �  B����    E�C��    �  ̐���    E�C��    �  V���2   E�C)�$     h���U    E�CF�E�A�    $   ,  ����U    E�CF�E�A�    4   T  ��L   E�CM�����-�B�B�B�B�A�      �  ֖��7    E�C       $   �  ���w    E�CG��d�B�A�(   �  <���{    E�CI���d�B�B�A�      �����    E�C�� $      ����   E�CE���A�       H  ����    E�Cx�     $   l  @���\    E�CF�L�A�       �  t���5   E�C,�   �  ����_    E�CV� ,   �  Ȟ���   E�CG����B�A�       $     ����P    E�CF�@�A�    $   ,  ����Z    E�CF�J�A�    $   T  ݠ��^    E�CF�N�A�       |  ���4    E�Ck�     �  '���v   E�Cm�$   �  }����    E�CF���A�       �  ����    E�C�� $     ݣ���    E�CF���A�       ,  J���*    E�Ca�     L  T���'    E�C^�     l  [���/    E�Cf�     �  j���;    E�Cr�     �  ����;    E�Cr�     �  ����:    E�Cq�     �  ����'    E�C^�       ����9    E�Cp�     ,  ڤ��9    E�Cp�     L  ���<    E�Cs�     l  ���=    E�Ct�     �  ,���>    E�Cu�     �  J���n    E�Ce�    �  ����;    E�Cr�     �  ����9    E�Cp�       ̥��9    E�Cp�     ,  ���9    E�Cp�     L  ����D    E�C{�     l  "���9    E�Cp�     �  ;���9    E�Cp�     �  T���9    E�Cp�     �  m���9    E�Cp�  $   �  ����a    E�CF�Q�A�          ����2    E�Ci�     4   Ѧ��T    E�CF�   P   	���X    E�CF�$   l   E����    E�CG����B�A�   �   ����T    E�CF�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    GCC: (Ubuntu 9.3.0-17ubuntu1~20.04) 9.3.0                                        �                    �                    �                 h  �                 �  �                 @" �                  0 �                                     ��                     ��_ cole _             ��                )        �           &         �           0    ��                7    ��                ?     #  �   �      G      � �           M      � �           S      � �           Y      � �           _      
 �           e       �           k      ' �           q      6 �           w      8 �           }      j �           �      x �           �      � �           �      � �           �      � �           �    ��                �      � �           �      � �           �      � �           �      � �           �    ��                �    ��                �    ��                �    ��                �      � �           �        �           �       �           �    ��                �    ��                �    ��                �    ��                �      8 �           �      T �           �      x �           c   ��                �     @" �          �      � �           �       �              ��                	   ��                �      4 �              ��                   ��                "   ��                +   ��                8   ��                A   ��                J   ��                S   ��                \   ��                f   ��                o   ��                x   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �    H" �          �   ��                �   ��                �   ��                �   ��                �   ��                �      8 �              ��                   ��                   ��                    ��                �      ` �           (   ��                0   ��                9   ��                C   ��                K   ��                B   ��                J   ��                R   ��                Z   ��                b   ��                j   ��                s   ��                |   ��                �   ��                �   ��                �   ��                �   ��                �    )�  �   �       �      x �           �   ��                �   ��                �    ��  �   �       �      p �           �      w �           �   ��                �   ��                �   ��                �    `" �          �   ��                [   ��                �   ��                �   ��                �      p �           �   ��                �   ��                �    T�  �   e       >    ��  �   �           [�  �   �      �    `" �              ��  �   =      	    `# �          �    ��  �   �       �   ��                �   ��                   ��                   ��                &   ��                �      x �           0   ��                9    `$ �   `       A   ��                �      � �           J   ��                Q   ��                Y   ��                b   ��                k   ��                r   ��                ~   ��                }   ��                |   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �      � �           �   ��                �    �$ �          �    �$ �          �    �  �   {       �    ��  �   �       �    =�  �   �      �   ��                �      � �           �   ��                �      � �           �      � �           �      � �           �   ��                �    A�  �   _       �      � �           �      � �           �      � �           �      � �           �   ��                   ��                   ��                   ��                   ��                $   ��                +   ��                ,   ��                3   ��                T   ��                ;   ��                D   ��                P   ��                [   ��                c   ��                �      � �           j   ��                p   ��                w   ��                �        �           ~   ��                �       �           �   ��                �       �           �   ��                �       �           x   ��                �        �              ��                �      ( �           �   ��                �      0 �           �   ��                �      8 �           �   ��                �      @ �           �   ��                �   ��                �      H �           �      Y �           �   ��                �      m �           �      ~ �                ��                �    h  �           �    P�  �   T       �    c  �         �    p�  �   \       �    �:  �   �       �    :�  �   {       �    
�  �   9           </  �   Z           h�  �   ;           ��  �   �           �a  �   �       (    "M  �   �       3    @% �          ,    �  �   7          r�  �   �       5    �$ �          <    *�  �   �      E    x"  �   �       O    B+  �   Z       W    "�  �   �       ^      �           f    ~.  �   �       �    <6  �   �       n    �$  �   �       r      �           w    ��  �   P       �    ��  �   �       �    �. �          �    �  �   �       �    ��  �   �       �    �$ �          �    D�  �   �      �    ��  �   U       �    �F  �   u       �    ��  �   w       �    =�  �   9       �    �. �          �    �  �   9       �    5�  �   ^       �    ` �          �    /�  �   �       4    B�  �   �       �    K�  �   [      �    t  �   :      �    Nv  �   �           �+  �   �       [
    �  �   �           H% �               R%  �   z      &    1�  �   w       -    �  �   �      7    LC  �   �       F    ?J  �   �      N    �  �   L       U    ��  �   v      �    ��  �   �       \    J�  �   U       d    ��  �   \       k    ��  �   Y       p    '�  �   M       w    �  �   K       
    �$ �          ~    �& �          �    �C  �   �      �    C�  �   <       �    ��  �   �       �    �  �   L      �    k�  �   G      �    �$ �          �    �R  �         �    `% �          �    �f  �   ]      �    �6  �   �       �    w�  �   K              �               �7  �   �          ]G  �   �           0 �               0Q  �   Z      )    �  �   �       /    &)  �   Z       8     ]  �   A       ?    b�  �   �       K    �M  �   2      R    n[  �   �       Z    >�  �   2      a    �$ �          �
    s�  �   �       f    iU  �   �       n    ��  �   �       v    ��  �   �       {    t�  �   O       �    �  �   5      �    A]  �   i       �    ��  �   P           Ӷ  �   �       �    �)  �   @       �    "\  �   �       �    ŗ  �   z       �    *e  �   �      �    �*  �   �       7     ` �           �    ��  �   �       �    ��  �   Y       �    \�  �   9       �    �(  �   Z       �    �/  �   h           �w  �   �          ��  �   �      �    ��  �   9           �$ �                 �          P
    @" �               �. �          %       �           ,     % �          5     ` �           ;    ��  �   �       B    �a  �   9       L    �^  �   g       
    N�  �   D       �	    ��  �   '       Z    ��  �   >       `    	�  �   T       g    -.  �   Q       o    ��  �   V       w    *�  �   �           9,  �   h      �    �]  �   U       �    '5  �         �    ��  �   n       �    ��  �   }       �    �4  �   �       �    
�  �   �       �    ��  �   9       �    �& �          �    �  �   S       �    \9  �   j      �    H�  �   k       �    Qi  �         Q
    @" �            	    S�  �   W       	    N  �   H      	    ��  �   �       	    �/  �   Z       "	    g�  �   �       )	    ��  �   �       5	    Nu  �          @	    �  �          K	    ]�  �   X       U	    �Z  �   �       \	    "w  �   �       m	    J�  �   ]       s	    ` �          z	    �l  �   D      �	    �. �          �	    `  �   �      �	    B�  �   �       �	    ��  �   �       �	       �           �	    ��  �   9       �	    5�  �   ;       �	    ��  �   b       �	    % �          �	    <"  �   <       �	    M�  �   K       �	    z�  �   *       �	    ,�  �   K       �	    ��  �   �       3    ��  �   /       �	    PV  �   r       �	    `*  �   @       �	       �           
    % �          :    ��  �   �       �    v�  �   a       
    C�  �         �
    §  �   S       
    !C  �   +       �    �X  �   �      k    2  �         $
    PT  �   �       ,
    ��  �   l       "    �V  �         6
    ��  �   �       V
    ��  �   9       =
    �F  �   I       C
    ��  �   e      O
    @" �           U
    ��  �   9       Z
     �  �   K       =    ��  �         `
    �;  �         o
    ��  �   Z       v
    ��  �   6      ~
    �  �   9       �
    =�  �   �       �
    ��  �   2       5    -�  �   �       �
    % �          �
    �{  �   i      �
    ,�  �   �       �
    �S  �   �       �
    �  �   '          ��  �   �       �	       �           �
    `& �          �
     % �          �
    ��  �   S       �
    �T  �   p       �
    �)  �   �       �
    �-  �   2       �
      �   @      �
    N   �           �
    �  �   C          p�  �   :           ��  �   u          ��  �   �           X0  �   '      #    ��  �   ]       *    (% �          6     ` �           3    <�  �   \      ;    O�  �   L       B    a�  �   Y       �       �           J    �  �   �       �
    f�  �   7       T    �-  �   Z       ]    0% �          d    ��  �   a       n    p�  �   U       �    �A  �         s    ��  �   �       ,    ]=  �   �      |    T^  �   i       �    ��  �   ;       �    �  �   3      �    `   �   �      �    �<  �   �       �    �  �   L       �       �           �    ��  �   U       �    �B  �   9       �    $_  �   �       �    ��  �   '       �       �           �    �b  �   ^           b�  �   �       �    ��  �   4       �    ?�  �   a       �    ��  �   �       �    ��  �   9       �    ��  �   +          �  �   =           ��  �   �          '�  �   r           �]  �   U       +    ��  �   L       0    ʏ  �   O       lib/setup.asm HEADER_MAGIC HEADER_FLAGS header crt0.c shell.c cmd_run .LC35 .LC36 .LC37 .LC38 .LC39 .LC40 .LC41 .LC42 .LC43 .LC44 .LC45 .LC46 .LC47 .LC48 dir.c .LC0 .LC1 .LC2 .LC3 gui.c font8x16.c window.c bmp.c font.c border.c file.c cfs.c alloc_spin_lock pipe.c path.c memcmp.c memcpy.c memset.c strcasecmp.c strcat.c strchr.c strcmp.c strcpy.c strcspn.c string.c strlen.c strncasecmp.c strncmp.c strncpy.c strpbrk.c strrchr.c strsep.c strspn.c strtok.c last.1481 strstr.c strdup.c memmove.c strcoll.c strerror.c ctype.c tolower.c toupper.c stdio.c fopen.c fclose.c fflush.c fputc.c fgetc.c fgets.c fputs.c fread.c fwrite.c remove.c rewind.c fseek.c feof.c ftell.c vfprintf.c vf vsprintf.c vsnprintf.c sn_buf putchar.c sscanf.c perror.c vfscanf.c character _buf.1638 fvalue _buf.1650 ungetc.c getchar.c freopen.c tmpnam.c _tmpnam rename.c itoa.c i2hex.c malloc.c calloc.c free.c realloc.c lldiv.c strtol.c atoi.c atol.c strtoul.c exit.c getenv.c qsort.c qscmp qses qsexc qstexc qs1 system.c strtod.c ftoa.c _precision atof.c strtof.c strtold.c abs.c ltoa.c utoa.c srand.c errno.c gmtime.c localtime.c strftime.c clock.c math.c pow.c sqrt.c atan.c acos.c asin.c floor.c ceil.c exp.c locale.c signal.c setjmp.c _GLOBAL_OFFSET_TABLE_ longjmp read_directory_blk drawstring strcpy log cmd_date sqrt setjmp clean_blk_enter put strtok_r stdout vsprintf wait_exit cmd_mov ungetc pwd_ptr cmd_del set_argv strerror utoa_r __m_i memmove __tm __realloc_r atol __window_puts getenv ceil errno floor strtold _infinity qsort fgets file_update file_read_block cmd_info call_loader shell memcpy cmd_table __window_clear BitMAP2 perror ltoa_r tolower system feof malloc remove fs_directory __window_putchar ldexp vsnprintf strtoul itoa __pipe__ stdgetc_r argv_pointer update_directory_entry _drawline fflush argc drawrect BitMAP eh_frame stdputc_r upath cmd_time tell_r strncasecmp border write_r strtol user flush_r strrchr utoa calloc strtod rewind_r atof cmd_shutdown seek_r strcat read_directory_entry cmd_new debug_o fseek __free_block_r cmd_version cmd_clear open_dir ftoa stdin font8x16 __m_c _start obj_list __end strstr write_blk get_file_name atan2 signal cmd_dir strcoll strncmp cmd_help write_sector draw_char_transparent pow strncpy put_pixel strcasecmp log10 _BLK_ realloc drawchar path_count open_file_r strtok remove_blk memcmp cmd_copy sscanf getfilename file_close pipe_write sigaction read_r file_write_block fread _ctype open_file addr search_blk_null strdup fopen sysgettmpnam localtime memset pwd main ftell srand fclose getchar close_r cmd_reboot __data ptr_mouse2 __free_r update_window getkeyw _vsputs_r strcmp color remove_file __bss atan fgetc drawchar_trans strtof strcspn asin ltoa setlocale stderr create_file strsep getkey __malloc_r _v_ mouse fputc open_r cmd_rename cmd_exit A__ call_function getpathname strftime i2hex lldiv cmd_cd fwrite __window vfscanf rewind freopen pipe_read cmd_echo pipe_r __block_r atoi __heap_r assert_fn gmtime strspn ctr0 drawstring_trans strlen __code toupper wcl filename_cmp clock read_super_block abs strchr fputs acos strchrnul frexp vfprintf strpbrk read_sector free setpath  .symtab .strtab .shstrtab .text .data .got .got.plt .data.rel.local .bss .eh_frame .comment                                                                                    �           �                             !                �                                          '                �          h                              ,             h  �   h                                   5             �  �   �      �                              E             @" �   0"     �                             J              0 �    0      0                             T      0                `     *                                                   0`     �,      
   �                 	                       �     8                                                   8�     ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ELF          >       �   @       0�         @ 8  @                   �      �    �       �                             �      �   `"       0                   0      0 �    0 �                          Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��  ���_ cole _          �      �            P �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           I��H�P% �   L�H�0% �   H�H�   �   L�H�  �   L�#H�  �   L�+�   �����H��H��H��H��L�������UH��AWSH��@��H�����I���      L�H�}�H�u�H�U�H�M�L�E�L�M�H���������H�H�U�H�H��     H�E�H�H�E�H��     H�H��     H�H� H��H��     H�H��     H�H��H��     H�H��     H�H�@H��H��     H�H�E�H��     H�H�E�H��     H�H�E�H��     H�H��     H�H��H��     H�I�߸    H�!e������H���H��     H�    H���������H�H� H��H��     H�H���������H�H� H��H���������H�H� H�։�I��H��������H��ЉE�E��I��H��������H��АH��@[A_]���UH��AWSH���   ��H�����I��      L�H�� ����    �    H��I��H�4u������H����E�    H��H���H��I��H���������H���H�E�H�Eȋ@H�       H�H�H��H�Eȋ@H�       H�H�H��H�� ���H���������H�43H��I�߸    I�5�������I�A��H���������H�H� H�E�H�E�H   � �? �    H��I��H�4u������H���H�E��PH�E��PH�E��PH�E��PH�E��@     H�E��@    H�E��PH�E��P(H�E��PH�E��P$H�E��@0    H�E��@,    H�E��@H   H�E��@L   H�E��@P    H�E��@T��� H���������H�H��H�E�H�PXH�E��@��H�E��@��H�E��@��H�E��@ ��H�E�I��A��� �I��H��������H���H�E��@��H�E��@��$��H�E��@ ��H�E�I��A���� �$   I��H��������H���H�E��@ ���E�H�E��@��"�E��E�    �E�   H�E��P �E�Ѓ��E�H�E��@��"�E��E�    �E�   H�E��P �E�E�Ѓ��E�H�E��@��"�E��E�    �E�   �    I��H���������H���H�E��    I��H���������H���H�E��    I��H���������H���H��x����   I��H���������H���H��p���H���������H�4H���������H�<I��H�"�������H���H��h���H��h��� ��   H��h����   �    H��I��H�'�������H���H��h���H��I��H�ً������H��Љ�d���H��h���H��I��H�ۊ������H��Ћ�d���H��h���H�E��   H��I��H�։������H���H�M��U��u�H�E�I�ȹ��� H��I��H��%������H���H��h���H��I��H���������H����%H���������H�<I�߸    H���������H���H���������H�4H���������H�<I��H�"�������H���H��h���H��h��� ��   H��h����   �    H��I��H�'�������H���H��h���H��I��H�ً������H��Љ�`���H��h���H��I��H�ۊ������H��Ћ�`���H��h���H�E��   H��I��H�։������H���H�M��U��u�H�E�I�ȹ��� H��I��H��%������H���H��h���H��I��H���������H����%H���������H�<I�߸    H���������H���H���������H�4H���������H�<I��H�"�������H���H��h���H��h��� ��   H��h����   �    H��I��H�'�������H���H��h���H��I��H�ً������H��Љ�\���H��h���H��I��H�ۊ������H��Ћ�\���H��h���H��x����   H��I��H�։������H���H�M��U��u�H��x���I�ȹ��� H��I��H��%������H���H��h���H��I��H���������H����%H���������H�<I�߸    H���������H���H�E�H��I��H�t!������H��п�   I��H���������H���H��P����E�    �E�    �E�    �E�    H�E�    �H���������H�H� �@������  ��H���������H�H� �@����u�E�H���������H�H� � 9E��l  H���������H�H� �@9E��O  H���������H�H� � �M��U��9��,  H���������H�H� �@�M��U��9��  �}���   H�M��U��u�H�E�I�ȹ    H��I��H��%������H��Ѓ}� ucH�E�H��P���H���������H�4H��I��H��w������H���H���������H�H� �   H��P���H�uй   I���rH�EЉE���   �E�   ���rH�M��U��u�H�E�I�ȹ��� H��I��H��%������H���H�M��U��u�H��x���I�ȹ��� H��I��H��%������H���H���������H�H� � 9E��l  H���������H�H� �@9E��O  H���������H�H� � �M��U��9��,  H���������H�H� �@�M��U��9��  �}���   H�M��U��u�H�E�I�ȹ    H��I��H��%������H��Ѓ}� ucH�E�H��P���H���������H�4H��I��H��w������H���H���������H�H� �   H��P���H�uй   I���rH�EЉE���   �E�   ���rH�M��U��u�H�E�I�ȹ��� H��I��H��%������H���H�M��U��u�H��x���I�ȹ��� H��I��H��%������H���H���������H�H� � 9E��l  H���������H�H� �@9E��O  H���������H�H� � �M��U��9��,  H���������H�H� �@�M��U��9��  �}���   H�M��U��u�H��x���I�ȹ    H��I��H��%������H��Ѓ}� ucH�E�H��P���H���������H�4H��I��H��w������H���H���������H�H� �   H��P���H�uй   I���rH�EЉE���   �Eܹ   ���rH�M��U��u�H�E�I�ȹ��� H��I��H��%������H���H�M��U��u�H�E�I�ȹ��� H��I��H��%������H����E�    H�Eȋ@9E���   H�Eȋ@�E�H�Eȋ@H�       H�H�H��H�Eȋ@H�       H�H�H��H�� ���H���������H�43H��I�߸    I�5�������I�A��H�U�H�� ���H��H��I��H�m ������H�����u�����UH��AWSH��P��H�����I�1�      L�H�}�H���������H�H� H�Eؿ  � I��H���������H���H�E��E�    �E�    H�E�H�E�H�E�H��������H�4H��I��H�"�������H���H��     H�H��     H�H��u*H��������H�<I�߸    H���������H����0  H��     H��   �    H��I��H�'�������H���H��     H�H��I��H�ً������H��ЉE�H��     H��    �    H��I��H�'�������H���H��     H��U�H�Eо   H��I��H�։������H��ЋU�9�t*H� �������H�<I�߸    H���������H����P  H�E�H�.�������H�4H��I��H�߀������H���H�E�H�E�H��H�1�������H�<I�߸    H���������H���H�.�������H�4�    I��H�߀������H���H�E�H�E��
   �    H��I��H���������H��ЉE�H�.�������H�4�    I��H�߀������H���H�E�H�E��
   �    H��I��H���������H��ЉE�H�.�������H�4�    I��H�߀������H���H�E�H�E��
   �    H��I��H���������H��ЉE�H�E�H��I��H��z������H��Љ�H�PH�E�H�H�E�H�u�M��UȋE�I����H�8�������H�<I�߸    I���������I�A���E�    �   �E�    �yH�E�H�PH�U�� �E�H�E�H�PH�U�� �E�H�E�H�PH�U�� �E��E� H�E�H��   H�E��H�E؋P�E�Hc��E�H�I��H��I��H�������H��ЃE��E�9E��{����E��E�9E��b���H��     H�H��I��H���������H���H�E�H��I��H�O�������H��и    H��P[A_]���UH��H��0��H�����I���      L�H�}�H�u��U܉M�L�E�H���������H�H� H�E��E�H9E�}?H�E��@��H9E�}0H�E�H�E��E�H�E�H��H�E�H�H��    H�E�HE؉������UH��SH��@��H�����I�@�      Lۉ}ԉuЉỦM�L�E�L�M�f�E�  H�E�H�@H�E�H�E��@�E�}�u�E�    �E�    �   f�E� H�E��@�EȉE��H�H� H�E�H�� f�E�H�E�� ���E��J�E�f#E�f��t5�UЋE��Hc��UԋE��H�H�}��M�U�I��H��H�������H���f�e�m��}� y��E�H�E��@9E��b�����H��@[]���UH��AWSH��0��H�����I�)�      Lۉ}܉u؉UԉM�D�E�L�M��E�    �X�E�    �CH�E�L��   �M�H�E��P�u؋E��Hc��}܋E��H�H��I��H�������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I�z�      Lۉ}܉u؉UԉM�D�E�L�M��E�    �p�E�    �[H�E�H��   �E��E�i��E��A��H�E��P�M؋E��Hc��M܋E��H�I��D��H��I��H�������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I���      Lۉ}܉u؉UԉM�D�E�L�M��}� �[  �}� �Q  �E�    �>H�E�L��   �M�H�E��P�E�Hc��}܋E��H�H��I��H�������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E����Hc��}܋E��H�H��I��H�������H��ЃE��E�;E�|��E�    �AH�E�H��   �M�H�E��P�u؋E��Hc��E�H�I��H��I��H�������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E��Hc��}܋E����H�H��I��H�������H��ЃE��E�;E�|���H��0[A_]���UH��AWSH��@��H�����I�	�      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}��  �E�    ��   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��   �E�f#E�f��tDH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�������H����BH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�������H���f�e�m��}� �[����E�H�E��@9E��	�����H��@[A_]���UH��SH��8��H�����I���      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H��������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I���      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}���   �E�    �   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��W�E�f#E�f��tBH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�������H���f�e�m��}� y��E�H�E��@9E��T�����H��@[A_]���UH��SH��8��H�����I���      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H�������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I��      L�H�}ȉuĉU��M�D�E�D�M�H���������H�H� H�E�H�E�H   � �? �    H��I��H�4u������H����E�    �U�H�E��P4�UH�E��P8�UH�E��P<H�E��@H   H�E��@L   H�E��P<H�E��PP�UH�E��PTH���������H�H��H�E�H�PXH�E��@D    H�E��PDH�E��P@�U�H�E��P�U�H�E��P�U�H�E��P �U�H�E��P�U H�E��P`�} u�E�   H�E��@�P�H�E��P(H�E��P�E�)ЍP�H�E��P$H�E��@0   �E����H�E��P,H�E��@��H�E��@��H�E�I���Ѻ    �    I��H��,������H���H�E��@4��H�E��@����H�E�I��A�ȹ   �   �   H��������H��Ѓ}� u:H�E��@����H�E�I��A���� �   �   �   H��������H����8H�E��@����H�E�I��A���� �   �   �   H��������H��Ѓ}� t}H�E��@����H�U��E�I��A���� ����   �   H��������H���H�E��@4��H�E��@���ƋE��H�U�I��A�ȹ   ��ƿ   H��������H���H�E��@8A��H�E��@$��H�E��@(��H�E��@,��H�E��@0��H�E�I��H��������H���H�E�H��I��H��z������H������E�H�E�H�pHH�E��@��E܉������)Љ�H�E�H���u�I��A���� ������   ��H��H�-������H���H��H�E��@����H�E�I��A�    �   �   �   H�>������H���H�E�H�PHH�E��@��H���u�I��A���� ������   �ƿX   H�������H���H��H�E�H�PHH�E��@��(H���u�I��A���� ������   �ƿ-   H�������H���H��H�E�H�e�[A_]���UH��AWSH��0��H�����I���      L�H�}�H�u�H�E��P0H�E��@Ѓ�P�E�H�E��P,H�E��@Ѓ��E��E�P   �E�   �E�    �E���� H�E�H��I��H��z������H��ЉE�H�E�L�@H�M؋U܋E���������p��E�<�E��������ƋE���)ƋE��H�E�H���u�M��A�ȉщ�H��H�R������H���H���H�e�[A_]���UH��H����H�����I���      L�H�}��   H�E�H���r�����UH��H����H�����I�G�      L�H�}������UH��H����H�����I��      L�H�}�H�U��BD    H�U��JDH�U��J@H�U��R8A��H�U��R$��H�U��R(A��H�U��R,��H�U��R0��H�U�I��D��I��������J��А����UH��SH��(��L�����I���      Mډ�f�E�H���������I�H� H�E�H���������I�H��H�E�H�PXH�E�@(�P�H�E�@H���к    ��E�H�E�@$�P�H�E�@L���к    ��E�H�E�P<H�E�PPH�E�PD�E�9�rH�E��@D    H�E�@@�PH�E�P@H�E�P@�E�9�r9H�E��@D    H�E�PDH�E�P@H�E�H��H��!������I����E��  f�}���   H�E�@D����   H�E�@D�P�H�E�PDH�E�H�xHH�E�pTH�E�@PH�U�J,H�U�RLA��H�U�R@A��ʃ���H�U�J0H�U�RHA��H�U�RDA��ʃ�A��H���u�I��A������D�޿    H��������I���H����   f�}�	uH�E�@D�PH�E�PD��   f�}�
u!H�E��@D    H�E�@@�PH�E�P@�   f�}���   H�E�H�xHH�E�pTH�E�PPH�E�H,H�E�@LA��H�E�@@A��ȃ���H�E�H0H�E�@HA��H�E�@DA��ȃ�A���E�H���u�I��A���щ�D�މ�H��������I���H��H�E�@D�PH�E�PD�E�H�]�����UH��H����H�����I���      L؉}�H���������H�H� H�E��U�H�E��P<�����UH��SH��(��H�����I��      L�H�}�H�}� t=H�E�H�E��&H�E�H�PH�U�� f�����H�e"������H���H�E�� ��u���H��([]���UH��AWSH��P��H�����I��      L�H�}��u��U��M�L�E�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H�W�������H�<I�߸    H���������H��Ҹ�����6  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H�e�������H�<I�߸    H���������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�}�������H�<I�߸    H���������H��Ҹ   ��   �E�    �   �E�    �   �}� tNH�E�H��   H�E��P�M��E���E��Hc��M��E���E��H��M�I��H��I��H�������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�������H��ЃE��}� �U����E��}� �;����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��P��H�����I�&�      L�H�}��u��U��M�D�E�L�M�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H�W�������H�<I�߸    H���������H��Ҹ�����3  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H�e�������H�<I�߸    H���������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�}�������H�<I�߸    H���������H��Ҹ   ��   �E�    �   �E�    �   �}� tKH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�������H��ЃE��}� �X����E��}� �>����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��0��H�����I�C�      Lۉ}܉u؉U�H�M��E�    �   �E�    �t�U�������E��H���������H�Hڋ��E�}� tBH�E�H��   H�EȋP�MԋE��Hc��M؋E��H��M�I��H��I��H�������H��ЃE��}�~��E��}��o�����H��0[A_]���UH��AWSH��@��H�����I�g�      Lۉ}̉uȉUĉM�L�E��E���� �E�``` �E���� �EĉE��ẺE܋E��E؋EȉEԋE؍P��E��xH�M��E�I��A�    �   ��I��H�>������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H�>������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H�>������H��ЋEԍP��E܍pH�M��E�I��A�    �Ѻ   ��I��H�>������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H�>������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H�>������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H�>������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H�>������H��ЋEԍP��E܍p�M��E�ȃ�H�M�I��A�    �Ѻ   ��I��H�>������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H�>������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H�>������H��ЋE؍P��M܋E�ȍp��E���H�M�I��A�    �   ��I��H�>������H��АH��@[A_]���UH��AWSH����H�����I�5�      Lۉ}�H�u�H�E�� ��H�E��@9�sH�E��P#H�E��@9�r"H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@��u)H���������H�H��E�H�։�H��/������H���H�E�H�PH�E��@#��H�H�E�H�PH�E�H�@�U�H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  H�E��@��u0H���������H�H� H��t�E�����I��H�e"������H��ЋE�H��[A_]���UH��H����H�����I���      L�H�}��E�    H�E�@��u]H�E�@'�PH�E�P'��H�E�P#H�E�@'9�r�H�E�H�PH�E�@'��H��H�H�E�H�PH�E�H�@� ���E��   H�E�@��tH�E�@��uiH�E�@#��u������ZH�E�P'H�E�@#9�r������AH�E�H�PH�E�@'��H�H�E�H�PH�E�H�@� ���E�H�E�@'�PH�E�P'�E�����UH��H����H�����I���      L�H���������H�H� H�E��E�    H�E��@��uWH�E��P#H�E��@'9�w�    �AH�E�H�PH�E��@'��H�H�E�H�PH�E�H�@� ���E�H�E��@'�PH�E��P'�E�����UH��H����H�����I��      L�H���������H�H� H�E��E�    H�E��@��uXH�E��@'�PH�E��P'��H�E��P#H�E��@'9�r�H�E�H�PH�E��@'��H��H�H�E�H�PH�E�H�@� ���E��E�����UH��AWH��(��H�����I�m�      L�H�}�H�u�H�U����u�    �(H�M�H�U�H��H��I��H�\K������H���H�E�H�E�H��(A_]���UH��AWSH�� ��H�����I���      L�H�}�H�}� u
������   H�}� tH�E؋@����tH�E��@"<t������zH�E؋@%�   ��u�    �cH�E؋@#H�U؋J�    ��E�H�E؋@��@��u�U�H�E؉�H��I��H��U������H���H�E�H��I��H��R������H��ЉE�E�H�� [A_]���UH��AWSH����H�����I��      L�H�}�H�}� u������0H�E�H��H��3������H���H�E�H��I��H��S������H���H��[A_]���UH��AWSH�� ��H�����I���      Lۉ}�H�u�H�}� u
�������  H�EЋ@��u
�    �  H�EЋ@��tH�EЋ@��tH�EЋ@��u!H�UЋE�H�։�H��/������H����y  H�EЋ@����unH�EЋP#H�EЋ�+  9�wYH�EЋ�+  ��tKH�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��E�U�H�EЉ�H��I��H��T������H����H�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U܈H�E�� ��H�EЋ@��9�r3H�EЋ@����H�EЉPH�E�f�   H�E�H��H��3������H���H�EЋ@#�PH�EЉP#H�EЋP#H�EЋ�+  9�vH�EЋ�+  �PH�EЉ�+  H�EЋ@���H�EЉP�    H�� [A_]���UH��AWH��(��H�����I���      L�H�}�H�}� u
������  H�E؋@��u
�    �v  H�E؋@��tH�E؋@��tH�E؋@��u"H�E�H��H�1������H��ЉE�E��0  H�E؋P#H�E؋�+  9�r
������  H�E؋@����ulH�E؋P#H�E؋�+  9�wWH�E؋�+  ��tIH�E؋@����H�E؉PH�E؋@#H�U؋r�    ���E�U�H�E؉�H��I��H��T������H���H�E؋@#H�U؋J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@� ���E�H�E�� ��H�E؋@��9�rH�E؋@����H�E؉PH�E�f�   H�E؋@#�PH�E؉P#�E�H��(A_]���UH��SH��H��H�����I���      L�H�}ȉuĉU�H�M�H�}� u�    �y�E�    H�E�H�E��E�    �FH�E�H��H�j7������H��ЉE؃}��u�E�    �u��4H�E�H�PH�U��U؈�E��E��E��E��E�9�w��E�    �u�H��H[]���UH��SH��H��H�����I���      L�H�}ȉuĉU�H�M�H�}� u�    �l�E�    H�E�H�E��E�    �9H�E�H�PH�U�� ���E�H�U��E�H�։�H�N5������H��ЃE��E��E��E��E�9�w��E�    �u�H��H[]���UH��H����H�����I�F�      L�H�}�H�u��U�}�tZ�}�|�}� t�}�t�nH�E���H�E��P#H�E���H�E��P'�RH�E��@#H�U��H�E��P#H�E��@'H�U��H�E��P'�(H�E���+  H�U�)Љ�H�E��P#H�E��P#H�E��P'�H�E��@#H�U��J�    ��Љ�H�E�f��    ����UH��H����H�����I�h�      L�H�}�H�}� u�    �	H�E��@#������UH��H����H�����I�'�      L�H�}�H�}� t7H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@����H�E��P������UH��H��(��H�����I���      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H��(��H�����I�i�      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H����H�����I��      L�H�}��E�_   �(�E�Hc�H�E�H�� < u�E�Hc�H�E�H��  �m��}� y����    ����UH��H����H�����I���      L�H�}�H�E�H�E�H�E�H�E��H�E�� </uH�E�H��H�E�H�E�H�E�� ��u�H�E�����UH��H��0  ��H�����I�A�      L�H������H������H������H�E�H������H�E�H������H�E��E�    �?H�E�� ��u�E�Hc�H�E�H��  �H�E�H�PH�U��U�Hc�H�U�H�� ��E��}�_~��E�    �-H�E�H�PH�U��H�E�H�PH�U�� 8�t�   ��E��}�_~͸    ����UH��SH�� ��H�����I�\�      L�H�}�H�u�H�E؋PH�E؋@ЉE�E�H�U����H�     H�H�¾   H�6<������H��ЉE�}� t
�������   �E�    ��   �E�%�  ��H�     ��H؋���uf�E�%�  ��H�     ��H��������E�H�U����H�     H�H�¾   H��<������H��ЉE�}� t������r�E��m�E�%�  =�  uE�E��E�H�U����H�     H�H�¾   H�6<������H��ЉE�}� t�������E�H�E؋@$9E����������H�� []���UH��H����H�����I�ӿ      L؉}��u�H�U�H�M�    ����UH��AWSH��0��H�����I���      Lۉ}�H�u�H�U�H�EȋPH�Eȋ@ЉE�H�Eȋ@ �E܉E�ЉE�   �    H�     H�<I��H�4u������H����E�    �B�U�E�Љ�H�EЋ ��H�     H��   H��<������H��ЉE��}� u�E�H�EȋP �E�9�w���H��0[A_]���UH��H����H�����I���      L�H�}�H�u�H�U��R��H�U����H�U�H��H��   I�6<������J� ������UH��AWSH��`��H�����I�P�      L�H�}�H�u�H�U�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�E�H�E�H�E�H��I��H��r������H��ЉE�H�E��@,�E��9  H�E�H�E��H�E�� </uH�E��  H�E��H�E�H�E�� ��u׋U�H�E��@ H�M��	��H�M���H�6<������H��ЉE؃}� t#H�E�H��I��H�O�������H��и    ��   �E�    �f�E���Hc�H�E�H�H�E�H�E��@a��t5H�E��@b����@��t#H�E�H�U�H��H��H��=������H��ЉE���E������}� t�E��}�?~����}� u+�}�?%H�EЋ@k�E�H�E��@ �E؉E�ЉE�m��	�E�    �
�}� �����H�E�H��I��H�O�������H��ЋE�H��`[A_]���UH��AWSH��P��H�����I�;�      L�H�}�H�u�H�U��M�L�E�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�Eغ    �    H��I��H�4u������H��ЋU�H�E��@ H�M��	��H�M؉�H�6<������H��ЉE�}� t#H�E�H��I��H�O�������H��и������   �E�    �T�E���Hc�H�E�H�H�E�H�E��@a��t#H�E�H�U�H��H��H��=������H��ЉE���E������}� t�E��}�?~����}� u:�}�?4�E���Hc�H�E�H�H�EȺ�   H��H��I��H��t������H�����E�����H�E�H��I��H�O�������H��ЋE�H��P[A_]���UH��AWSH��P��H�����I�q�      L�H�}�H�u�H�U�H�E���C  ��u
������	  H�E���C  ��@v/H���������H�<I�߸    H���������H��Ҹ������  H�E��PH�E��@ЉE�H�E���?  H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�Eغ    �    H��I��H�4u������H��ЋU�H�E��@ H�M��	��H�M؉�H�6<������H��ЉEԃ}� t!H�E�H��I��H�O�������H��ЋE��  H�E���C  ��H��H��H�E�H�H�E�H�EȺ`   �    H��I��H�4u������H���H�E�H��+H��H�I=������H���H��H�E�H��H��I��H��w������H����E�    �"H�UȋE�H����uH�UȋE�H�� �E��}�_~�H�E��@` H�E���+  H�EȉPo�U�H�E��@ H�M��	��H�M؉�H��<������H��ЉE�H�E�H��I��H�O�������H��ЋE�H��P[A_]���UH��AWSH��`��H�����I��      L�H�}�H�u�H�U��S  I��H���������H���H�E�H�EкS  �    H��I��H�4u������H���H�E��PH�E��@ ��H�EЉP�    I��H���������H���H�U�H�BH�E��PoH�EЉ�+  H�E��PH�EЉ�/  H�E��P H�EЉ�3  H�E��H�EЉ�G  �    I��H���������H���H�U�H��K  H�E�H��K  �    �    H��I��H�4u������H���H�E��@k�E�    I��H���������H���H�E��E������E�    �E�    ��  �   I��H���������H���H�U�H��K  �M�Hc�H��H�H�H�E�H��K  �U�Hc�H��H�H� H�E�H�E��   �    H��I��H�4u������H����E�    �<  H�E��@ �E��H�E��@�H�E��P�E�H�H�4�    H�E�H�ʉH�EЋ�;  �PH�EЉ�;  �E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E�;E�ts�E�H�U����H�U�H��H�¾   H�6<������H��ЉE��}� t:H�E�H��I��H�O�������H���H�E�H��H��S������H��и    �   �E��E�H�E��@�����E�    ��U�E�H��    H�E�HЋ �E�}��u	�E�������E��}��  ������}��t�E��}��  � �����H�E�H��I��H�O�������H���H�E�H��`[A_]���UH��AWSH��p  ��H�����I���      L�H������H�������   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H������H�E�H��H��I��H��p������H���H�U�H�E�H��H��I��H�?s������H��п�   I��H���������H���H��     H�H��     H���   �    H��I��H�4u������H��п   I��H���������H���H�E�H�EȺ   �    H��I��H�4u������H���H�E�H�E�H�E��   �    H��I��H�4u������H����E�    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ ���    Hǅ���    Hǅ���    Hǅ���    Hǅ ���    Hǅ(���    Hǅ0���    Hǅ8���    Hǅ@���    HǅH���    HǅP���    HǅX���    Hǅ`���    Hǅh���    Hǅp���    Hǅx���    H�E�    H�E�    H������H������H��H��I��H��w������H���������<wt������<au�E�   H�E��@   H�E��     H�U�H�E�H��H��H�CA������H��ЉE�}� t_H��     H�H��I��H�O�������H���H�E�H��I��H�O�������H���H�E�H��I��H�O�������H��и    �  H�E�H�U�H�M�H�E�H��H��H��A������H��ЉE��}� u_H��     H�H��I��H�O�������H���H�E�H��I��H�O�������H���H�E�H��I��H�O�������H��и    �  H�EȋU��P,H��     H�H�M�H�U�H�u�I�ȹ    H��H��C������H��ЉE�}����   �}� tqH��     H�H������H�U�H�u�A�    H��H�qZ������H���H��     H�H������H�U�H�u�I�ȹ    H��H��C������H��ЉE�}� ��   H��     H�H��I��H�O�������H���H�E�H��I��H�O�������H���H�E�H��I��H�O�������H��и    ��  �}� t_H�E�H��I��H�O�������H���H��     H�H��I��H�O�������H���H�E�H��I��H�O�������H��и    �r  H��     H�H�U�H�M�H��H��H��G������H���H�E�H�}� ��   H��     H�H��H�E�H��+�`   H��H��I��H��t������H���H�E�H��+H��H��<������H���������<wt������<+t������<au
H�E��@"�H�E��@"H�E��@   H�EȋP,H�E���?  H��     H��PsH�E���C  ������<auH��     H��PoH�E��P#H�E�H��I��H�O�������H���H��     H�H��I��H�O�������H���H�E�H��I��H�O�������H���H�E�H��p  [A_]���UH��AWSH��@��H�����I�Q�      L�H�}��   I��H���������H���H�E�H�E�   �    H��I��H�4u������H���H�E�H�E�H�E�   �    H��I��H�4u������H���H�E��@   H�E��     H�U�H�E�H��H��H�CA������H��ЉE܃}� t H�E�H��I��H�O�������H��и�����AH�U�H�M�H�E�H��H��H��E������H��ЉE�H�E�H��I��H�O�������H��ЋE�H��@[A_]���UH��AWSH�� ��H�����I��      L�H�}�H�E�H�@H��I��H�O�������H����E�    �TH�E�H��K  �U�Hc�H��H�H� H��t?H�E�H��K  �U�Hc�H��H�H� H��I��H�O�������H��ЃE��}��  ~���H�E�H��K  H��I��H�O�������H���H�E�H��I��H�O�������H���H�E�    �    H�� [A_]���UH��H�� ��L�����I��      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H�6<������I� ������UH��H�� ��L�����I�F�      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H��<������I� ������UH��AWSH��   ��H�����I�l�      L�H��x���H��p�����l����   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H��x���H�E�H��H��I��H��p������H���H�U�H�E�H��H��I��H�?s������H��п   I��H���������H���H�E�H�EȺ   �    H��I��H�4u������H���H�E�H�E�H�E��   �    H��I��H�4u������H���H�E��@   H�E��     H�U�H�E�H��H��H�CA������H��ЉE��}� t_H��     H�H��I��H�O�������H���H�E�H��I��H�O�������H���H�E�H��I��H�O�������H��и�����-  H�E�H�U�H�M�H�E�H��H��H��A������H��ЉE��}� u_H��     H�H��I��H�O�������H���H�E�H��I��H�O�������H���H�E�H��I��H�O�������H��и�����  H�EȋU��P,H�EȋPH�Eȋ@ЉE�H�EȋP,H�Eȋ@ �ЋE�ЉE��    I��H���������H���H�E�H�E��    �    H��I��H�4u������H��ЋU�H�Eȋ@ H�M��	��H�M���H�6<������H��ЉE��E�    �E�    �   �E���Hc�H�E�H�H�E��E�;�l���}~H�E��@a��ta�E���Hc�H��p���H�H�E���   H��H��I��H��t������H��ЋE���Hc�H��p���H�H��H��<������H��ЃE����E��}�?�e�����H�E�H��I��H�O�������H���H�E�H��I��H�O�������H���H�E�H��I��H�O�������H��ЋE�H�Đ   [A_]���UH��AWSH��`��H�����I���      L�H�}�H�u�H�U�H�M�D�E�H�E�H�E�H�Eغ�   �    H��I��H�4u������H���H�E�H��H�I=������H���H��H�E�H��H��I��H��w������H����E�    �"H�U؋E�H����uH�U؋E�H�� �E��}�_~�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉEп    I��H���������H���H�E�H�EȺ    �    H��I��H�4u������H��ЋU�H�E��@ H�M��	��H�Mȉ�H�6<������H��ЉEă}� t!H�E�H��I��H�O�������H��ЋE���  �E�    �$�E���Hc�H�E�H�H�E�H�E��@a��t�E��}�?~���H�E��@a���G  �}�?�=  �U�H�E؉PsH�E��@a��E���H�E؈PbH�U�H�E�H��H��H��>������H���H�U؉BkH�E؋@k���uOH�E�H��H���������H�<I�߸    H���������H���H�E�H��I��H�O�������H��и   ��   �E���@��t$H�E؋@kH�U�H�M�H�Ή�H�Z@������H���H�M�H�E຀   H��H��I��H��t������H��ЋU�H�E��@ H�M��	��H�Mȉ�H��<������H��ЉEĐH�E�H��I��H�O�������H��и    �JH�E�H��I��H�O�������H���H�E�H��H���������H�<I�߸    H���������H��Ҹ����H��`[A_]���UH��AWSH��P��H�����I��      Lۉ}�H�u�H�U��    I��H���������H���H�E��E�    �E��E��E������E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E��E܋E�;E���   �}� tV�E�H�U����H�U�H��H�¾   H��<������H��ЉẼ}� t#H�E�H��I��H�O�������H��и�����?  �E�H�U����H�U�H��H�¾   H�6<������H��ЉẼ}� t#H�E�H��I��H�O�������H��и������   �E��E�E��E��E�   H�E��@�����E�    ��U�E�EȋE�H��    H�E�HЋ �E�E�H��    H�E�H��     �}��uL�E�H�U����H�U�H��H�¾   H��<������H��ЉE̐H�E�H��I��H�O�������H��ЋE��6�E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��Y���H��P[A_]���UH��AWSH��   ��H�����I�̟      L�H��h����   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H��h���H�E�H��H��I��H��p������H���H�U�H�E�H��H��I��H�?s������H��п   I��H���������H���H�E�H�E��   �    H��I��H�4u������H���H��p���H�E�H�E��   �    H��I��H�4u������H���H�E��@   H�E��     H�U�H�E�H��H��H�CA������H��ЉE�}� t<H�E�H��I��H�O�������H���H�E�H��I��H�O�������H��и    ��  H�E�H�U�H�M�H�E�H��H��H��A������H��ЉE��}� u<H�E�H��I��H�O�������H���H�E�H��I��H�O�������H��и�����d  H�E��U��P,H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE��    I��H���������H���H�E�H�E��    �    H��I��H�4u������H��ЋU�H�E��@ H�M��	��H�M���H�6<������H��ЉE�}� tSH�E�H��I��H�O�������H���H�E�H��I��H�O�������H���H�E�H��I��H�O�������H��ЋE��l  �E�    �   �E������E���Hc�H�E�H�H�E�H�E��@a��t!H�E�H�U�H��H��H��=������H��ЉE�}� u9H�E��@a �U�H�E��@ H�M��	��H�M���H��<������H��ЉE�}� ��E��}�?�k����}� tPH�E�H��I��H�O�������H���H�E�H��I��H�O�������H���H�E�H��I��H�O�������H��ЋE��uH�E��@kH�U�H�M�H�Ή�H��]������H��ЉE�H�E�H��I��H�O�������H���H�E�H��I��H�O�������H���H�E�H��I��H�O�������H��ЋE�H�Đ   [A_]���UH��H����H�5����I�m�      Lމ}�E�E��}� u�E��   �E����rH�(     H�H�(     H�����UH��H����H�����I��      L�H�}��   H�E�H���r�����UH��AWH����H�����I�њ      L�H�     H�H�U�H�      H�    H��      �    H�M�   �    H��I��H�4u������H��ѐH��A_]���UH��AWSH��P��H�����I�I�      Lۉ}��u��}� u
�    ��  H�      H�H=�   v%H�0�������H�<I�߸    H���������H��ҐH��      ���u�H��      ��PH��      ��E����E�E�%�  ��t�E��E�    �E�    �E�    �}� t�E��   �E�   �K  �}��  �=  H�     H�H�E�H�E�    �E�    �  H�E؋@����   H�E؋@9E���   H�E�H�H�E؋@��H�H�E�H�E؋@+E���H�E؉PH�E؋P�E��H�E؉PH�E�H�E�H�     H�H�E��E�    �mH�E؋@��tH�E��E��WH�E�H�E�H�E�H�E�H�E�H�@H�PH�E�H�PH�E��@   H�E�H�U�H�H�E��U��PH�E�H�U�H�P�E���!�}��   ~��H�E��E��}��   ������E�   ���}� ��   H�     H�H�E��E�    �~H�E؋@��tH�E��E��hH�E�H�E��E��H��d������H���H�E�H�E�H�U�H��E��E���H�E��PH�E��U��P�E���+E���H�E��PH�E�H�@   ��}��   �u���H��      �    H�      H�H�PH�      H�H�E�H��P[A_]���UH��SH��(��H�����I�$�      L�H�}�H�}� ��  �H��      ���u�H��      ��PH��      �H�E�H�E�H�     H�H�E��E�    �M  H�E�H� H9E�tH�E��E��2  H�E�H�E�H�      H�H�P�H�      H�H�E؋@��uH�E�H��H��d������H����   H�E؋@��uH�E�H�@H�E�H�E�H�@H�P�H�E�H�PH�E�H�@H��tH�E؋@����   H�E�H�@H��uRH�E�H� H��H��d������H���H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    ��}��   �������H��      �    ��H��([]���UH��AWH��H��L�����I�"�      M�H�}��u�H�E�    �E�    H�}� u�E��   ��H��e������I� ���8  �H��      A� ��u�H��      A� �PH��      A� H�     I� H�E�H�E�H�E��E�    �   H�E�H� H9E�t
H�E��   H�E�H�E��E�   H�E��P�E��=   v@H�      I� �U�H�E�H��H�h�������I�< M�Ǹ    I���������M�A����H�E�H� H�E�H�E��P�E��H�E��P�E��}��   �X���H��      A�     �}� u�E��   ��H��e������I� ���H�E�H��HA_]���UH��H�� ��H�����I���      L�H�}�H�u��E�    H�E�H�E��   H�E�� ��H�E��@9�sH�E��P#H�E��@9�rH�E��@#    H�E�f�   H�E�H�PH�E��@#��H�H�E�H�PH�E�H�PH�U�H�U�H�R� �H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  �E��}��E����E�����UH��H�� ��H�����I���      L�H�}�H�u��E�    H�E�H�E�H�E��@'�PH�E��P'H�E��P'H�E��@9�rH�E��@'   �H�E��P#H�E��@'9�r�H�E��@'�P�H�E��P'�JH�E�H�PH�E��@'��H�H�E�H�PH�E�H�PH�E�H�HH�M���H�E��@'�PH�E��P'�E��}�~��E�����UH��AWSH��0��H�����I���      L�H�}�H���������H�H� H�E�H�E�H�E�H�E�H��I��H��z������H��ЉE�H�E�H��I��H��z������H��ЉE؋U܋E��=   ~
������   H�E�� </uH�E��E�H�HE�H�m�H�E�� </tH�E�H�E�H�PH�U�� /�H�E�H�U�H�E�H��H��I��H��w������H���H�E�H��I��H��z������H��Љ�HE�H�m�H�E�� </u	H�E��  �H�E�H�E��  �    H��0[A_]���UH��AWSH����H�����I�L�      L�H���������H�H� H��I��H��z������H��Ѓ�w
�    �   H���������H�H� H�E�H�E�H��I��H��z������H��Љ�HE��H�E�H�P�H�U��  H�E�� </u�H���������H�H� H��I��H��z������H��Ѓ�vH�E��  �    H��[A_]���UH��AWSH��0��H�����I�`�      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
�    ��  H�E�H��I��H��z������H��ЉE�E�H�H�P�H�E�H�� </u�E�H�H�P�H�E�H��  �}� 
�    �  �}���   H�E�H��� <:u%H�U�H�E�H��H��I��H��w������H����K  H���������H�<I��H�)�������H���H��H�E�H��H��I��H��w������H���H�E�H��I��H��z������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H��w������H����   H���������H�<I��H�)�������H���H��H�E�H��H��I��H��w������H���H�E�H��I��H��z������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H��w������H���H�E�H��0[A_]���UH��H����H�����I� �      L�H�}�H�E�H�E�H�}� u�    �+�E�    �H�E�� </u�E�H�E�H�E�� ��u�E�����UH��AWSH��0��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
������   H�E�H��I��H��z������H��ЉE�E�H�HE�H�m��H�E�� </tH�m�H�E�� ��t�E�P��U�����H�E�H�U�H�E�H��H��I��H��w������H���H�E��  �    H��0[A_]���UH��H��8��H�����I�͋      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �CH�E�H�PH�U�� ���E�H�E�H�PH�U�� ���E�E�+E�E�}� u�}� t
�m��}� u��E�����UH��H��8��H�����I�7�      L�H�}�H�uЉŰẺE�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M����E��P��U���u�H�E�����UH��H�� ��H�����I���      L�H�}���U��E�E��E�H�E�H�E��H�E�H�PH�U��U��m��}� u�H�E�����UH��AWSH��0��H�����I�[�      L�H�}�H�u�H�E�H�E�H�E�H�E��E�    H�E�H�PH�U�� ����I��H�փ������H��ЉE�H�E�H�PH�U�� ����I��H�փ������H��ЉEԋE�+EԉE܃}� u�}� t뗋E�H��0[A_]���UH��AWSH����H�����I���      L�H�}�H�u�H�E�H��I��H��z������H��Љ�H�E�H�H�E�H��H��I��H��w������H���H�E�H��[A_]���UH��H�� ��H�����I�)�      L�H�}�u�H�E�H�E��H�E�� ��9E�uH�E��H�E�H�E�� ��u۸    ����UH��H�� ��H�����I�Ȉ      L�H�}�H�u�H�E�H�E�H�E�H�E��3H�E��H�E�� 8�u!H�E�� ��H�E�� ��Ѕ�u�    �'H�E�H�PH�U��H�E�H�PH�U�� 8�t����������UH��H��0��H�����I�.�      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E��  H�E�����UH��AWH��(��H�����I���      L�H�}؉uԋU��҉Uԃ}� uOH�U�H��I��H��z������H��҉�H�E�H���   H�E�� ��tH�E�� ��9E�u	H�E��   H�E�H�E؃�H��űE�i��E�H�E�H�E��H�E�H�E� ������H�E� ��!�%������u%H�E� 3E䍐����H�E� 3E���!�%������t�H�E�H�E��H�E�H�E�� ��tH�E�� ��9E�u�H�E�H��(A_]���UH��H��@��H�����I���      L�H�}�H�u�H�U�H�U�H�U������   H�U�H�������   H�E�    H�E�    H�E�    H�E�    �H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�t�H�E�H+E��'H�U����H�Uȉ�H��H�Ax������H���H+E�����UH��H����H�����I�R�      L�H�}�H�E�H�E��H�E�H�E�� ��u�H�E�H+E�����UH��AWSH��@��H�����I��      L�H�}�H�u��U�H�E�H�E�H�E�H�E��E�    �kH�E�H�PH�U�� ����I��H�փ������H��ЉE�H�E�H�PH�U�� ����I��H�փ������H��ЉEԋE�+EԉE܃}� u�}� t
�m��}� u��E�H��@[A_]���UH��H��(��H�����I�>�      L�H�}�H�u��U�H�E�H�E�H�E�H�E��}� u)������2H�E�H�PH�U��H�E�H�PH�U�� 8�u�m��}� u����E�����UH��H��8��H�����I���      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �!H�U�H�BH�E�H�E�H�HH�M����E��E�9E�w�H�E��  �E�����UH��AWH����H�����I�?�      L�H�}�H�u�H�M�H�U�H��H��I��H�ly������H��҉�HE�H�E�� ��tH�E���    H��A_]���UH��AWH��(��H�����I�͂      L�H�}؉u�H�U�H��I��H��z������H��҉E��U�H�E�H�H�E��E�    �H�E�� ��9E�uH�E��H�m��E��E�9E�wڸ    H��(A_]���UH��H��0��H�����I�<�      L�H�}�H�u�H�E�H� H�E�H�}� u�    �vH�E�H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u,�}� u
H�E�    �H�E�H���  H�E�H�U�H�H�E���}� u������UH��H��@��H�����I��      L�H�}�H�u�H�E�H�E�H�E�    H�E�    H�E�    H�E�    H�E�� ��u
�    ��   H�E�H��� ��u+�H�E�H�E��H�E�� 8�t�H�E�H+E��   H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�u�H�E�H+E�����UH��H��8��H�����I�L�      L�H�}�H�u�H�U�H�}� uH�E�H� H�E�H�}� u
�    ��   �H�E�H�PH�U�� ���E�H�E�H�E��
�E�;E�u��H�E�H�PH�U�� ���E��}� uۃ}� uH�E�H�     �    �   H�E�H��H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u4�}� u
H�E�    �H�E�H��H�E�H�E��  H�E�H�U�H�H�E���}� u������UH��H����H�����I�      L�H�}�H�u�H�u�H�M�H�       H�H��H��������H�������UH��AWSH�� ��H�����I��~      L�H�}�H�u�H�E�H��I��H��z������H��ЉE��2�U�H�M�H�E�H��H��I��H�'t������H��Ѕ�uH�E��H�E�H�E�� ��uø    H�� [A_]���UH��AWSH�� ��H�����I�#~      L�H�}�H�E�H��I��H��z������H��Ѓ��E�E��I��H���������H���H�E�H�}� u�    �$�U�H�M�H�E�H��H��I��H��t������H��АH�� [A_]���UH��H��8��H�����I��}      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��U�H�E�H�H�E�H�E�H;E�v[H�E�H;E�sQH�E�H�E��E�HE��H�m�H�m�H�E��H�E��H�E�H;E�u��'H�U�H�BH�E�H�E�H�HH�M���H�E�H;E�u�H�E�����UH��AWH����H�����I��|      L�H�}�H�u�H�M�H�U�H��H��I��H�,w������H���H��A_]���UH��AWH����H�����I�l|      Lډ}�H���������H�<I�׸    H���������H�������UH��H����H�����I�|      L؉}��U���H���������H�Hc��������t�E� �E�����UH��H����H�����I��{      L؉}��U���H���������H�Hc��������t�m� �E�����UH��AWSH��0��H�����I�q{      L�H�}ȉuĉU��M��U�H�E�H��H���������H�<I�߸    I���������I�A��H�E�H��I��H���������H���H�E�H�E� �E�H�E� 9E�u��H��0[A_]���UH��AWSH�� ��H�����I��z      L�H�}�H�u�H�E�� ��u�    �LH�E�� <wuH�E�H��I��H���������H���H�U�H�E�H��H��I��H��3������H���H�E�H�E�H�� [A_]���UH��AWH����H�����I�:z      L�H�}�H�U�H��I��H��4������H���H��A_]���UH��AWH����H�����I��y      L�H�}�H�U�H��I��H��3������H���H��A_]���UH��AWH����H�����I��y      L؉}�H�u�H�M��U�H�Ή�I��H�N5������H���H��A_]���UH��AWSH�� ��H�����I�Py      L�H�}�H�}� u������VH�E�H��I��H�j7������H��ЉE�H�E؋@��u+H���������H�H��E�H�։�I��H�N5������H��ЋE�H�� [A_]���UH��AWH����H�����I��x      L؉}�H�u�H�M��U�H�Ή�I��H�N�������H���H��A_]���UH��AWH����H�����I�fx      L�H�}�H�U�H��I��H���������H���H��A_]���UH��AWSH��@��H�����I�x      L�H�}ȉu�H�U�H�}� u	H�E��  H�E�H�E�H�E�H�E��E�    H�E�H��I��H�j7������H��ЉEԃ}����   H�E��@��u7�}�u�}� ~+H���������H�H��E�H�։�I��H�N5������H��Ѓ}�
tk�E�;E�}E�}�u�}� ~H�E�H;E�vH�m��m��:�}��^���H�E�H�PH�U�UԈ�E��D����}�u�}� ~�m���E��)�������}�~	H�E��  ��Eԉ�H�E�H�E�H��@[A_]���UH��AWSH�� ��H�����I��v      L�H�}�H�u�H�}� u�    �^�E�    �2�E�Hc�H�E�H�� ��H�U�H�։�I��H�N�������H��ЃE�H�E�H��I��H��z������H��ЋU�9�w��E�H�� [A_]���UH��AWH��(��H�����I�v      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I�99������I�A��H��(A_]���UH��AWH��(��H�����I��u      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I��9������I�A��H��(A_]���UH��AWH����H�����I�bu      L�H�}�H�U�H��I��H�"`������H���H��A_]���UH��AWH����H�����I�u      L�H�}�H�U�H��I��H��;������H��ҐH��A_]���UH��AWH��(��H�����I��t      L�H�}�H�u��U܋U�H�u�H�M�H��I��H��:������H���H��(A_]���UH��H����H�����I�tt      L�H�}�H�}� u������!H�E��P#H�E���+  9�r�������    ����UH��AWH����H�����I�t      L�H�}�H�U�H��I��H��;������H���H��A_]���UH��AWSH��`  ��H�����I��s      L�H������H������H�������E�    �E�    �  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H���������H���	E�}���  �E�H��    H��h  H�H��h  H�>��H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E��E�H������H�։�I��H�9�������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�}� t(H������H�E�H��H��I��H�2�������H����O  H������H��H���������H�<I��H�2�������H����   H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E�H�������E�H�։�I��H���������H���H������H������H��H��I��H�2�������H����w  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������
   H��H��I��H�q�������H���H������H������H��H��I��H�2�������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������   H��H��I��H�>�������H���H������H������H��H��I��H�2�������H����  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�EȾ   H��fHn�I��H�,�������H���H������H������H��H��I��H�2�������H����]  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eк
   H��H��I��H���������H���H������H������H��H��I��H�2�������H����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ
   H��H��I��H�q�������H���H������H������H��H��I��H�2�������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ   H��H��I��H�q�������H���H������H������H��H��I��H�2�������H����G  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�E�   H��fHn�I��H�,�������H���H������H������H��H��I��H�2�������H����   H������H�ƿ%   I��H�9�������H��ЋE�Hc�H������H�� ��H������H�։�I��H�9�������H����4�E�Hc�H������H�� ��H������H�։�I��H�9�������H��ЃE��E�Hc�H������H�� ��������    H��`  [A_]���UH��H����H�����I�?k      L؉��E��E�    �E��S��%wa��H��    H��a  H�H��a  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��j      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H�$�������L��Љ�<�����<���H���   A_]���UH��H�� ��H�����I��i      L�H�}�H�u�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E�����UH��AWSH��  ��H�����I�8i      L�H������H������H��x����E�    H������H�E�f�E�  �E� �E�    �/  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H���������H���	E܃}���  �E�H��    H�`  H�H�`  H�>��H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E��E�H�U�H�E�H��H��H�J�������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H�}� t'H�U�H�E�H��H��H�J�������H���H�E��e  H�E�H���������H�4H��H�J�������H���H�E��7  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E�H�������E�H�։�I��H���������H���H������H�E�H��H��H�J�������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������
   H��H��I��H�q�������H���H������H�E�H��H��H�J�������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������   H��H��I��H�>�������H���H������H�E�H��H��H�J�������H���H�E��3  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�E��   H��fHn�I��H�,�������H���H������H�E�H��H��H�J�������H���H�E��x  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�E��
   H��H��I��H���������H���H������H�E�H��H��H�J�������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ
   H��H��I��H�q�������H���H������H�E�H��H��H�J�������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ   H��H��I��H�q�������H���H������H�E�H��H��H�J�������H���H�E��e  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�Eо   H��fHn�I��H�,�������H���H������H�E�H��H��H�J�������H���H�E��   H�E�H���������H�4H��H�J�������H���H�E�fǅ����  �E�Hc�H������H�� ������H������H�E�H��H��H�J�������H���H�E��8�E�Hc�H������H�� �E�H�U�H�E�H��H��H�J�������H���H�E��E��E�Hc�H������H�� �������H�E��  H�U�H������H)�H��H�Ā  [A_]���UH��H����H�����I�i`      L؉��E��E�    �E��S��%wa��H��    H��X  H�H��X  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��_      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H���������L��Љ�<�����<���Hc�H�����H��  ��<���H���   A_]���UH��AWH���   ��L�����I��^      M�H����������H�����H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H����������H�����H��M��H�#�������L��Љ�<�����<���H���   A_]���UH��AWSH��0��H�����I��]      L�H�}؉u�H�U�H�M��}�   v
�    �   H�U�H�E�H��H�      H�<I��H���������H��ЉE�}���  ~�   �I�E�E�}� ~:�U�H�E�H�      H�4H��I��H��t������H��ЋE�Hc�H�E�H��  �E�H��0[A_]���UH��AWH����H�����I��\      L؉}�H���������H�H�
�U�H�Ή�I��H�N�������H���H��A_]���UH��AWSH�� ��H�����I��\      L�H�}�H�}� tj�E�    �?H���������H�H��E�Hc�H�E�H�� ��H�։�I��H�N�������H��ЃE�H�E�H��I��H��z������H��ЋU�9�w���H�� [A_]���UH��AWH���   ��L�����I��[      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H�$�������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I��Z      M�H��8���H��0���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�H���������I�<M�׸    H���������L�������UH��AWH����H�����I�^Z      L�H�}�H�U�H��I��H�X�������H��ҐH��A_]���UH��AWH��(��H�����I�Z      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H�ׇ������H��Ѹ    H��(A_]���UH��AWH��(��H�����I��Y      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H�ׇ������H����H�E�H�E�� < tH�E�H   H9E�sH�E�� <
u�H�E��  H�E�H;E�����H��(A_]���UH��AWSH��0��H�����I�
Y      L�H�}�H�uЉỦM�H�     H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H�ׇ������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H�     H�H�E�H�     �0H�     �D �}�u-�U�H�E�    H��I��H���������H���H�U�H��   �}�u+�U�H�E�    H��I��H�ʹ������H��Љ�H�EЉ�[�}�u,�U�H�E�    H��I��H�ʹ������H��Љ�H�E�f��)�U�H�E�    H��I��H�ʹ������H��Љ�H�EЈ�    H��0[A_]���UH��AWSH��0��H�����I�fW      L�H�}�H�uЉỦM�H�     H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H�ׇ������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H�     H�H�E�H�     �0H�     �D �}�u'H�E�H��I��H��������H����Z�H�E�� �+�}�u%H�E�H��I��H��������H���fH~�H�U�H��    H��0[A_]���UH��SH��8��H�����I�+V      L�H�}�H�u�H�U��E�    �E�    ��  �E�    �E�Hc�H�E�H�� ������%��  �E��E�Hc�H�E�H�� ������lu�E��E�   �E�Hc�H�E�H�� ����H�$�������H���	E�}��o  �E�H��    H�@O  H�H�5O  H�>��H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H��������H�����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H�E�������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H����?  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��������H�����   H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��������H����jH�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H������E��E�Hc�H�E�H�� ��������E�H��8[]���UH��H����H�����I��Q      L؉��E��E�    �E��S��%wa��H��    H�/L  H�H�$L  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I�!Q      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H�ȩ������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I�6P      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H�ȩ������L��Љ�<�����<���H���   A_]���UH��H����H�����I�FO      L؉}�H�u�H�}� u������w�}��u������jH�E��@#��tH�E��@#�P�H�E��P#H�E��@#H�U��J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U���E�����UH��AWSH����H�����I��N      L�H���������H�H� H��I��H�j7������H��ЉE�}��t+H���������H�H��E�H�։�I��H�N5������H��ЋE�H��[A_]���UH��AWH��(��H�����I�N      L�H�}�H�u�H�U�H���������H�<I�ϸ    H���������H�������UH��H����H�����I��M      L�H�}��	   H�E�H���r�����UH��SH����H�����I�tM      L�H�}�H�}� u.H�     H�<H�F�������H���H�     H��H�E�H��H�F�������H���H�E�H��[]���UH��AWSH��0��H�����I��L      L�H�}�H�u�H�E�H���������H�4H��I��H�"�������H���H�E�H�}� u
������   �E�    H�E�H��I��H��z������H��ЉE܃}�`~	�E�   �$H�E�H�P+H�E�H��H��I��H��w������H���H�E��@���H�E��PH�E�H��I��H���������H��ЋE�H��0[A_]���UH��H��0��H�����I��K      L؉}�H�u�H�E�H�E��E܉E��E�    �}� y,H�E�H�PH�U�� -�}�   �u�E�����E���E��؉E�H�E�H�E�M�Hc�Hi�gfffH�� ��������)�����)��ʉЍH0H�E�H�PH�U�ʈ�E�Hc�Hi�gfffH�� ����)ЉE�}� u��}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWSH��@��H�����I��J      L�H�}�H�u��U�H�}� u#H�E�H�E�H�E�H�PH�U�� 0H�E��  �  H�E�H�E؋E�Hc�H�E�H�H�E��3H�E؃��E�H�m��}�	~�7   ��0   �U��H�m���H�E�H�E�H;E�wËE�Hc�H�E�H��  H�E�H�E��E�    �8H�E�� <0uH�E��"H�U�H�E�H��H��I��H��w������H�����E��E�;E�|�H�E�H�E�H�E�H��I��H��z������H��Љ�H�E؋E�H�U�)Љ�H�M�H�E�HȾ    H��I��H�4u������H���H��@[A_]���UH��AWH����H�����I�?I      L؉}�U�    ��I��H��e������H���H��A_]���UH��AWH����H�����I��H      L؉}�u�U��U��I��H���������H���H��A_]���UH��AWH����H�����I��H      L�H�}�H�U�H��I��H��h������H��ҐH��A_]���UH��AWH����H�����I�WH      L�H�}�u�M�H�U��H��I��H��j������H���H��A_]���UH��H����H�����I�H      L؉}�u�E��}�E��E��}�ЉE��}� x�E���y�E����E��E�+E�E��!�}� y�E���~�E����E��U��E�ЉE�H�E�����UH��H�� ��H�����I�~G      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H�� ��H�����I��F      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H��H��H�����I�*F      L�H�}�H�u��U�H�E�H�E�H�E�H�PH�U�� ���E�E���H���������H�H������ ��uǃ}�-u�E�   H�E�H�PH�U�� ���E��"�E�    �}�+uH�E�H�PH�U�� ���E�}� t�}�u9�}�0u3H�E�� <xtH�E�� <XuH�E�H��� ���E�H�E��E�   �}� u�}�0u�   ��
   �E��}� t	H��   ������H�E�E�Hc�H�E�H�H��H�ЉE؋E�Hc�H�E�H�H��H�E�}� t�}� ~�E�)E�H�E��]�H�E�    �E�    �E���H���������H�H��������t�m�0�[�E���H���������H�H���������5  �E���H���������H�H��������t�7   ��W   )E�E�;E���   �}� ��   �}� tgH�E�H;E�|H�E�H;E�u0�E�;E�~(�E�����H�E�   �H���������H�� �����   �E�   �E�H�H�U�H��H�E��E�H�H)E��eH�E�H;E�H�E�H;E�u-�E�;E�~%�E�����H�E����H���������H�� �����$�E�   �E�H�H�U�H��H�E��E�H�HE���H�E�H�PH�U�� ���E��y������H�}� t�}� t
H�E�H���H�E�H�U�H�H�E�����UH��AWH����H�����I��B      L�H�}�H�M�
   �    H��I��H�ʹ������H���H��A_]���UH��AWH����H�����I��B      L�H�}�H�M�
   �    H��I��H�ʹ������H���H��A_]���UH��AWAVAUATSH����H�����I�EB      L�H�}�H�uȉU�L�eп    L��L�`� �؉���H���������H�H������ ��uЃ�-u�   L��L�`� �����+uL��L�`� �؃}� t�}�u-��0u(A�$<xt	A�$<XuI�D$� ��I���E�   �}� u��0u�   ��
   �EċE�Hc������    H��I�ǋE�Hc������    H��H�Љ�A�    A�    ����H���������H�H��������t��0�T����H���������H�H��������tz����H���������H�H��������t�7   ��W   )�;]�}GE��x
M9�wM9�u��9�~A������A�   �E�H�L��Hc�I�L��L�`� ���;������E��yA�����H���������H�� "   �	����tI��H�}� tE��tI�D$��H�E�H�U�H�L��H��[A\A]A^A_]���UH��H����H�����I�@      L؉}��   �   ���r����UH��AWSH����H�����I��?      L�H�}�H�E�H���������H�4H��I��H�,w������H��Ѕ�uH���������H�H� ��    H��[A_]���UH��AUATSH�� ��H�����I�O?      L�H�}�H�u�H��     ��E�L�e�H�]�E�,$L��L�`��H��H�XD�(�m��}� uې�H�� [A\A]]���UH��H��8��H�����I��>      L�H�}�H�u�H�U�H��     ��E�H�E�H�E�H�E�H�E�H�E�H�E�H�E�� ���E�H�E�H�PH�U�H�U���H�E�H�PH�U�H�U���H�E�H�PH�U��U���m��}� u�������UH��SH��H��H�����I�*>      L�H�}�H�u�H��     ��E�H�E�H+E��EȋE�9E���  �E�����EȺ    ��E��EȋU�H�E�H�H�E�H�E�H�E�H�E�H�E�E�H�H��H��H�E�H�H�E�H�E�H;E�sjH�x     H�H�U�H�E�H��H���щEă}� u/�E�H�H��HE�H�U�H�E�H��H��H���������H�����  �}� y�E�H�HE���  �H�E�H;E���   H�x     H�H�U�H�E�H��H���щEă}� u)�E�H�HE�H�U�H�E�H��H��H���������H���뢃}� ��   H�E�H;E�uA�E�H�HE�H�U�H�M�H�E�H��H��H��������H��ЋE�H�HE�H�E�H�E��M���H�U�H�E�H��H��H���������H��ЋE�H�H��HE��E�H�HE���   �E�H�H��HE�����H�E�H;E���   H�E�H+E�H��H�E�H+E�H9�|4�E�Hc�H�E�H�H�E�H��H��H���������H���H�E�H�E������H�U�H�E�H��H��H���������H��ЋE�Hc�H�E�H�H�E������E�H�H��HE�H�U�H�M�H�E�H��H��H��������H��ЋE�H�H��HE�H�E�H�E������H��H[]���UH��H�� ��H�����I�9;      L�H�}��u�U�H�M�H�x     H�U�H��U�H��     ��U��U���H�U�H�H�U�H��H��H���������H��А����UH��AWH����H�����I��:      L�H�}�H���������H�<I�׸    H���������H��Ѹ����H��A_]���UH��H��@��H�����I�\:      L�H�}�H�u�H�U�H�U��H�E�H�U����H���������H�Hc���҃� ��u��E�    H�U���҃�+t��-u�E�   H�E�H����������E��E�    �E�    �E�    �;�M�H����������Y�H�U���҃�0�*��X��E�H�E��E�H�U����H���������H�Hc���҃���u�H�U����.uuH�E��?�M�H����������Y�H�U���҃�0�*��X��E�H�E��E��E�H�U����H���������H�Hc���҃���u��U�)U�}� uH��������f���  �}� t�E�H��������f(fW��E�H�U����etH�U����E��   �E�    H�E�H�U���҃�+t��-u�E�   H�E��E�    �%�M܉����҉�H�U���҃�0ʉU�H�E�H�U����H���������H�Hc���҃���u��}� t�U�)U���U�U�}����|	�}�   ~H�����������   H����������E��E�E܃}� yF�]��A�E܃���t&�}� y�E��^E��E���E��YE��E��}��E��Y��E��}� u�H�}� tH�E�H�U�H��E�����UH��H����H�����I�'7      L؉}�H�E�   �E�    �H�U�H��H��H�H�H�E��E��E�;E�|�H�E�����UH��AWSH��@��H�����I��6      L��E�H�}��u�H�}� u	H�E��  H�E�H�E�H�0�������f��f/E�v,H�E�H�PH�U�� -�E�H�8�������f(fW��E��E�H�H�������f/s�E��H,�H�E��/�E�H�H���������\��H,�H�E�H�       �H1E�H�E�H�E�H�E�H��x�H*��H��H���H	��H*��X��M��\�f(��EȋE���H���������H���H��x�H*��H��H���H	��H*��X��YE�H�H�������f/s�H,�H�E��*H�H���������\��H,�H�E�H�       �H1E�H�E�H�E�H�M�H�U�H�E�H�(�������H�43H��I�߸    I�5�������I�A��H�E�H��@[A_]���UH��AWH����H�����I��4      L�H�}�H�U�    H��I��H���������H���H��A_]���UH��AWH����H�����I��4      L�H�}�H�u�H�M�H�U�H��H��I��H���������H����Z�H��A_]���UH��AWH��(��H�����I�14      L�H�}�H�u�H�M�H�U�H��H��I��H���������H����E��E�H��(A_]���UH��H����H�����I��3      L؉}��E����3E�)�����UH��H��@��H�����I��3      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�    H�}� y>H�E�H�PH�U�� -H�       �H9E�uH��������H�E�H�E��H�E�H��H�E�H�E�H�E�H�M�H�gfffffffH��H��H��H��H��?H)�H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U��ʈH�M�H�gfffffffH��H��H��H��H��?H)�H��H�E�H�}� u�H�}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U߈H�E�H;E�w�H�E�����UH��AWH��8��H�����I�)2      L�H�}�H�uЉU�H�U�H�U�H�}� yH�U�H�JH�M��-H�]�H�U�H�U��}�u$H�M�H�u�   H��I��H�>�������H����H�M�H�U�H��H��H�S�������H���H�E�H��8A_]���UH��H��0��H�����I�|1      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E�H�M�H���������H��H��H��H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U�ʈH�E�H���������H��H��H��H�E�H�}� u�H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWH��8��H�����I��0      L�H�}�H�uЉU�H�U�H�U�H�U�H�U��}�u$H�u�H�M�   H��I��H�>�������H����H�M�H�U�H��H��H�x�������H���H�E�H��8A_]���UH��H����H�����I��/      L؉}������UH����H�����I��/      Lظ   ]���UH��H����H�����I��/      L�H�}��    ����UH��H����H�����I�n/      L�H�}�H���������H�H� ����UH��H����H�����I�3/      L�H�}�H���������H�H� ����UH��H�� ��H�����I��.      L�H�}��u�H�U�H�M�    ����UH����H�����I��.      Lظ    ]���UH��H����H�����I��.      L��E�H�P�������f������UH��H����H�����I�^.      L��E�H�P�������f������UH��H����H�����I�%.      L��E��}�H�P�������f������UH��H����H�����I��-      L��E�H�}�H�P�������f������UH��H����H�����I��-      L��E��M�H�P�������f������UH��H��(��H�����I�n-      L��E��M��E��U��U��E��E��E������������������������������]��E�����UH��H����H�����I� -      L��E����E����]��E�����UH��H����H�����I��,      L��E�H�X�������f������UH��H����H�����I��,      L��E�H�`�������f������UH��H����H�����I�S,      L��E�H�h�������f������UH��H����H�����I�,      L��E�H�p���������E��E�����UH��H����H�����I��+      L��E�H�x�������f������UH��H����H�����I��+      L��E�H���������f������UH��H����H�����I�d+      L��E�H���������f������UH��H����H�����I�++      L��E�H���������f������UH��AWH����H�����I��*      L��E��E�H���������H�f(�fHn�I��H���������H���H��A_]���UH��H����H�����I��*      L؉}�H�u�    ����UH��AWH����H�����I�]*      Lډ}�H�u�H���������H�<I�׸    H���������H�������UH��AWH��(��H�����I�	*      Lى}�H�u�H�U�H���������H�<I�ϸ    H���������H�������UH��AWSH�� ��H�����I��)      L�H�}�H���������H�<I�߸    H���������H����E�    �.�E�H�H��    H�E�HЋ ��I��H���������H��ЃE��}�?~̸����H�� [A_]���UH��AWH����H�����I�)      L�H�}�u�H���������H�<I�׸    H���������H�����f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f�                                                                    ~ � � � � � � � � ~             ~ � � � � � � � � ~                 l � � � � | 8                   8 | � | 8                   < < � � �   <                < ~ � � ~   <                      < <              � � � � � � � � � � � � � � � �           < f B B f <           � � � � � � � � � � � � � � � �        2 x � � � � x             < f f f f <  ~               ? 3 ? 0 0 0 0 p � �              c  c c c c g � � �               � < � < �             � � � � � � � � � � �               > � >                  < ~    ~ <                f f f f f f f   f f              � � � {                | � ` 8 l � � l 8  � |                       � � � �              < ~    ~ <  ~              < ~                           ~ <                      �                         0 ` � ` 0                         � � � �                       ( l � l (                      8 8 | | � �                   � � | | 8 8                                                 < < <                  f f f $                             l l � l l l � l l           | � � � |   � � |               � �   0 ` � �             8 l l 8 v � � � � v           0 0 0 `                             0 0 0 0 0 0               0         0                   f < � < f                         ~                                    0                     �                                                           0 ` � �             8 l � � � � � � l 8              8 x       ~             | �    0 ` � � �             | �   <    � |               < l � �                 � � � � �    � |             8 ` � � � � � � � |             � �     0 0 0 0             | � � � | � � � � |             | � � � ~     x                                                       0                  0 ` 0                      ~     ~                     ` 0      0 `             | � �                       | � � � � � � � |              8 l � � � � � � �             � f f f | f f f f �             < f � � � � � � f <             � l f f f f f f l �             � f b h x h ` b f �             � f b h x h ` ` ` �             < f � � � � � � f :             � � � � � � � � � �             <         <                   � � � x             � f f l x x l f f �             � ` ` ` ` ` ` b f �             � � � � � � � � � �             � � � � � � � � � �             | � � � � � � � � |             � f f f | ` ` ` ` �             | � � � � � � � � |           � f f f | l f f f �             | � � ` 8   � � |             ~ ~ Z       <             � � � � � � � � � |             � � � � � � � l 8              � � � � � � � � � l             � � l | 8 8 | l � �             f f f f <     <             � � �   0 ` � � �             < 0 0 0 0 0 0 0 0 <               � � � p 8                 <         <          8 l �                                                   �       0                                     x  | � � � v             � ` ` x l f f f f |                   | � � � � � |                < l � � � � v                   | � � � � � |              6 2 0 x 0 0 0 0 x                   v � � � � � |  � x       � ` ` l v f f f f �                 8      <                        f f <       � ` ` f l x x l f �             8         <                   � � � � � � �                   � f f f f f f                   | � � � � � |                   � f f f f f | ` ` �             v � � � � � |                � v f ` ` ` �                   | � ` 8  � |              0 0 � 0 0 0 0 6                    � � � � � � v                   � � � � � l 8                   � � � � � � l                   � l 8 8 8 l �                   � � � � � � ~   �             � �  0 ` � �                 p                                        p         p                       v �                        8 l � � � �                               ��� ��� ~~~                                 uuu ��� ��� ���                                 ��� ��� ��� ��� ;;;                          ��� ��� ~~~ ��� ���                         ��� ��� ���     ��� ���                         ��� ���      ��� ��� ppp                 @@@ ��� ���         III ��� ���                 ��� ��� ��� ��� ��� ��� ��� ���                 ��� ���                 zzz ��� ���         ``` ��� ���                     ��� ���         ��� ��� MMM                     ��� ��� bbb     ��� ���                         ||| ��� ���      ��C00 01 02 03 04 05 06 07 08 09 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 %s:%s r console.bmp open error
 folder.bmp edit.bmp term.bin  explore.bin  editor.bin       r error: fopen
 error: fread
 
  %s
    width %d height %d sig %d %lx
 BitMAP error
 Not suport BitMAP 4-bit Not suport BitMAP > 8-bit  Entrada maior que o limite
 Erro ao criar o arquivo "%s"
       Error ao criar o arquivo "%s", atingio o limite de arquivos na entrada de directorio
   Panic: __malloc, sem espaco na tabela de alocacao
      panic: realoc sem espaco, %lx size = %d %d
 PWD strerrorr
                      (((((�AAAAAABBBBBB                                �Dubug: %s %x %x
        (null)  "�������L�������З��������������6������������������������������"�������"�������"�������"�������"�������"�������"�������"�������"�������"�������"�������P����������������������f�������f���������������������������������������������������������������������������������������������������������������������������������������{�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������(null) %        Ʀ�������������~�������9����������������������=�������=�������Ʀ������Ʀ������Ʀ������Ʀ������Ʀ������Ʀ������Ʀ������Ʀ������Ʀ������Ʀ������Ʀ����������������������Z���������������������Z���������������������������������������u���������������������������������������������������������������������������������������Q�������c�����������������������~���������������c�������������������������������������������������������������������������������Z���������������l�����������������������u�������panic: sscanf()
        �������Ѱ������6�����������������������������s�������s������������������������������������������������������������������������������������߲������K�������������������������������������!�������!�������!�������!��������������!�������!�������!�������!�������!�������!�������!�������!�������!�������!����������������������!���������������������!���������������!�������!�������!�������!�������!�������!�������!�������!�������!��������������!���������������!�������!��������������panic: freopen()
 r+ PWD call system funtion error. 
                 $@       �        %lu.%lu                �              �C                                                                        �_�
�@panic: signal()
 panic: sigaction()
 panic: setjmp()  panic: longjmp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �$ �     �     �   �- �   �$ �   �- �      �   % �      �     �   (% �   @% �   H% �                           h �   k �   n �   q �   t �   w �   z �   } �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �   � �    �    �    �   
 �    �    �    �    �    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          zR x�  ,      @����   E�CG����B�A�          L   �����   E�CJ��  ,   l   ����]   E�CG��J�B�A�          �   ����    E�C�� $   �   [��   E�CE��A�   $   �   H���    E�CG����B�A�$     ����    E�CG����B�A�(   4  n���   E�CG����B�A�   (   `  ���j   E�CG��W�B�A�       �  *���    E�CE���� (   �  ���   E�CG���B�A�       �  �	���    E�CE���� (      M
���   E�CG��q�B�A�   $   ,  ���   E�CG����B�A�   T  ���9    E�Cp�     t  ���+    E�Cb�     �  ����    E�C��     �  ���   E�CE����   �  ���I    E�C@�     �  ���u    E�CE�f�A�(     1���   E�CG����B�A�   (   H  ����   E�CG����B�A�   $   t  ����    E�CG����B�A�,   �  R��2   E�CG���B�A�       (   �  T��Z   E�CG��G�B�A�      �  ���   E�C�     ����    E�C��    8  ���    E�C��     X  ���p    E�CF�`�A�$   |  ����    E�CG����B�A�$   �  � ��r    E�CG��_�B�A�(   �  � ��   E�CG��	�B�A�   $   �  �"���   E�CF���A�          }$���    E�CE���A�    D  %���    E�CE���A�   h  �%���    E�C��    �  h&��A    E�Cx�      �  �&��i    E�C`�        �  �&��U    E�CL�    �  '��U    E�CL�      8'��i    E�C`�    ,  �'��g    E�C^�    L  �'���    E�C�� $   l  �(���   E�CE�{�A�      �  �)��9    E�Cp�  $   �  
*���    E�CG����B�A�   �  �*��^    E�CU� (   �  	+��   E�CG���B�A�   (   (  �,���   E�CG����B�A�   (   T  �.��]   E�CG��J�B�A�   (   �  �0��   E�CG��l�B�A�   (   �  4��D   E�CJ��.�B�A�   (   �  ,;��:   E�CG��'�B�A�   $     :<��    E�CG����B�A�   ,  =���    E�C��    L  �=���    E�C�� (   l  z>���   E�CJ����B�A�   (   �  =B��i   E�CG��V�B�A�   (   �  zE��H   E�CG��5�B�A�   (   �  �G��e   E�CJ��O�B�A�      	  �K��a    E�CX�    <	  L��9    E�Cp�      \	  )L���    E�CF�w�A�(   �	  �L��'   E�CG���B�A�   $   �	  �O��   E�CE���A�   $   �	  `Q���   E�CF���A�      �	  �R��    E�C��    
  �S���    E�C�� (   <
  ~T��O   E�CG��<�B�A�   $   h
  �U���    E�CG����B�A�(   �
  eV��C   E�CG��0�B�A�      �
  |X��k    E�Cb� $   �
  �X���    E�CG����B�A�     �Y���    E�C��    $  �Y��w    E�Cn�    D  TZ��b    E�CY� $   d  �Z���    E�CG����B�A�$   �  )[��z    E�CG��g�B�A�   �  {[��a    E�CX�    �  �[���    E�C��    �  6\��{    E�Cr� $     �\��+   E�CF��A�      <  �]��6   E�C-�   \  �^��L    E�CC� $   |  �^���    E�CG����B�A�   �  v_���    E�Cw�    �  �_��}    E�Ct� $   �  3`��r    E�CF�b�A�    $     }`���    E�CF���A�       4  �`���    E�C��    T  �a��3   E�C*�   t  �b��7   E�C.�   �  �c��W    E�CN� $   �  �c���    E�CG����B�A�$   �  Vd���    E�CG����B�A�     �d���    E�C�� $   $  pe��V    E�CF�F�A�       L  �e��P    E�CF�       l  �e��U    E�CL�    �  f��U    E�CL� $   �  8f���    E�CG����B�A�$   �  �f���    E�CG����B�A�$   �   g��K    E�CF�{�A�     $   $  Cg��K    E�CF�{�A�     $   L  fg��S    E�CF�C�A�    $   t  �g���    E�CG����B�A�$   �  h��S    E�CF�C�A�    $   �  ,h��K    E�CF�{�A�     ,   �  Oh��[   E�CG��H�B�A�       $     zi���    E�CG����B�A�$   D  �i��]    E�CF�M�A�    $   l  +j��]    E�CF�M�A�    $   �  `j��K    E�CF�{�A�     $   �  �j��L    E�CF�|�A�     $   �  �j��Y    E�CF�I�A�         �j��Y    E�CP� $   ,  k��K    E�CF�{�A�     (   T  4k���   E�CJ��{�B�A�       �  �s���    E�C��     $   �  t���    E�CI���A�       �  �t��l    E�Cc� (   �  .u���   E�CJ����B�A�         �}���    E�C��     $   <  ]~��   E�CI���A�    $   d  6���    E�CI���A�    $   �  ����    E�CG����B�A�$   �  ����\    E�CF�L�A�    $   �  �����    E�CG����B�A�$     ^����    E�CI���A�       ,  +����    E�CI�    $   L  ����L    E�CF�|�A�         t  Ђ��e    E�CF�U�A�    �  ����    E�CF���A�(   �  �����   E�CG����B�A�   (   �  ���=   E�CG��*�B�A�   $     ���\   E�CE�M�A�      <  L����    E�C�� $   \  ֊���    E�CI���A�    $   �  �����    E�CI���A�       �  f����    E�C�� $   �  �����    E�CG��z�B�A�   �  ]���Y    E�CF�         ����9    E�Cp�  $   4  �����    E�CE�q�A�    $   \  ����    E�CG����B�A�   �  ׎��G   E�C>�,   �  ����u   E�CG��b�B�A�       $   �  C���M    E�CF�}�A�     $   �  h���O    E�CF��A�     $   $  ����L    E�CF�|�A�     $   L  ����S    E�CF�C�A�       t  ޑ���    E�C�    �  F����    E�C��    �  В���    E�C��    �  Z���2   E�C)�$   �  l���U    E�CF�E�A�    $     ����U    E�CF�E�A�    4   D  Ɩ��L   E�CM�����-�B�B�B�B�A�      |  ژ��7    E�C       $   �  ���w    E�CG��d�B�A�(   �  @���{    E�CI���d�B�B�A�   �  �����    E�C�� $     ����   E�CE���A�       8  ����    E�Cx�     $   \  D���\    E�CF�L�A�       �  x���5   E�C,�   �  ����_    E�CV� ,   �  ̠���   E�CG����B�A�       $   �  ����P    E�CF�@�A�    $     ����Z    E�CF�J�A�    $   D  ���^    E�CF�N�A�       l  ���4    E�Ck�     �  +���v   E�Cm�$   �  �����    E�CF���A�       �  ����    E�C�� $   �  ����    E�CF���A�         N���*    E�Ca�     <  X���'    E�C^�     \  _���/    E�Cf�     |  n���;    E�Cr�     �  ����;    E�Cr�     �  ����:    E�Cq�     �  ����'    E�C^�     �  Ŧ��9    E�Cp�       ަ��9    E�Cp�     <  ����<    E�Cs�     \  ���=    E�Ct�     |  0���>    E�Cu�     �  N���n    E�Ce�    �  ����;    E�Cr�     �  ����9    E�Cp�     �  Ч��9    E�Cp�       ���9    E�Cp�     <  ���D    E�C{�     \  &���9    E�Cp�     |  ?���9    E�Cp�     �  X���9    E�Cp�     �  q���9    E�Cp�  $   �  ����a    E�CF�Q�A�         è��2    E�Ci�     $  ը��T    E�CF�   @  ���X    E�CF�$   \  I����    E�CG����B�A�   �  ����T    E�CF�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    GCC: (Ubuntu 9.3.0-17ubuntu1~20.04) 9.3.0                                        �                    �                    �                 h  �                 �  �                 `" �                  0 �                                     ��                     ��_ cole _             ��                )        �           �         �           0    ��                7    ��                B       �           H      " �           N      $ �           T      0 �           Z      < �           `      G �           f      P �           l      Z �           r      g �           x    ��                �      x �           �      z �           �      � �           �      � �           �      � �           �      � �           �    ��                �    ��                �    ��                �    ��                �      � �           �      � �           �      � �           �    ��                �    ��                �    ��                �    ��                �        �           �       �           �      @ �           P   ��                �     `" �          �      � �           �      � �           �    ��                �    ��                �      � �           �    ��                   ��                   ��                   ��                %   ��                .   ��                7   ��                @   ��                I   ��                S   ��                \   ��                e   ��                s   ��                }   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �    h" �          �   ��                �   ��                �   ��                �   ��                �   ��                �        �           �   ��                �   ��                   ��                   ��                �        �              ��                   ��                &   ��                0   ��                8   ��                /   ��                7   ��                ?   ��                G   ��                O   ��                W   ��                `   ��                i   ��                r   ��                z   ��                �   ��                �   ��                �    �  �   �       �      8 �           �   ��                �   ��                �    �  �   �       �      0 �           �      7 �           �   ��                �   ��                �   ��                �    �" �          �   ��                H   ��                �   ��                �   ��                �      0 �           �   ��                �   ��                �    H�  �   e       �    ��  �   �       �    O�  �   �      �    �" �          �    ��  �   =      �    �# �          �    ��  �   �       �   ��                �   ��                    ��                	   ��                   ��                �      8 �              ��                &    �$ �   `       .   ��                �      J �           7   ��                >   ��                F   ��                O   ��                X   ��                _   ��                k   ��                j   ��                i   ��                q   ��                z   ��                �   ��                �   ��                �   ��                �   ��                �      M �           �   ��                �    �$ �          �    �$ �          �    �  �   {       �    ��  �   �       �    1�  �   �      �   ��                �      Q �           �   ��                �      p �           �      x �           �      � �           �   ��                �    5�  �   _       �      � �           �      � �           �      � �           �      � �           �   ��                �   ��                �   ��                   ��                
   ��                   ��                   ��                   ��                    ��                A   ��                (   ��                1   ��                =   ��                H   ��                P   ��                �      � �           W   ��                ]   ��                d   ��                �      � �           k   ��                �      � �           r   ��                �      � �           s   ��                �      � �           e   ��                �      � �           l   ��                �      � �           y   ��                �      � �           �   ��                �      � �           �   ��                �        �           �   ��                �   ��                �       �           �       �           �   ��                �      - �           �      > �                ��                �    h  �           �    D�  �   T       �    	b  �         5    d�  �   \       �    �9  �   �       �    .�  �   {       �    ��  �   9       �    \�  �   ;       �    ��  �   �       �    �`  �   �           L  �   �           �  �   7      2    f�  �   �           �$ �               �  �   �      )    �  �   �       0      �           �    05  �   �       8      �           =    �  �   P       F    ��  �   �       M    �- �          S    ֢  �   �       D    ��  �   �       [    �$ �          `    8�  �   �      l    ��  �   U       q    �E  �   u           ��  �   w       �    1�  �   9       _
    X% �          �    �- �          �    ��  �   9       �    )�  �   ^       �    ` �          �    #�  �   �       Z
    6�  �   �       �    ?�  �   [      �    s  �   :      �    Bu  �   �       �	    	�  �   �       �    %�  �   w       �    @B  �   �       �    3I  �   �      �    ��  �   L       �    ��  �   v      z    ��  �   �       �    >�  �   U           ��  �   \           �  �   Y           �  �   M           ��  �   K       K	     % �              `% �          ,    �B  �   �      =    7�  �   <       C    ��  �   �       �	    �  �   �      M    �  �   L      U    _�  �   G      Z    % �          c    ~Q  �         m    �e  �   ]      �    �5  �   �       �    k�  �   K       �       �           �    �6  �   �      �    QF  �   �      �     0 �           �    $P  �   Z      �    �  �   �       �    �[  �   A       �    V�  �   �       �    �L  �   2      �    bZ  �   �       �    2�  �   2      �    % �          �    g�  �   �       �    ]T  �   �            ��  �   �           ��  �   �           h�  �   O            �  �   5          5\  �   i       $    �  �   P       1    ǵ  �   �       )    [  �   �       0    ��  �   z       7    d  �   �      �     P �           L    �  �   �       T    ��  �   Y       Z    P�  �   9       i    �v  �   �      r    ��  �   �          ��  �   9       w    % �          }       �          �	    `" �           �    �- �          �       �           �     % �          �     P �           �    ��  �   �       �    �`  �   9       �    �]  �   g       �	    B�  �   D       $	    ��  �   '       �    ��  �   >       �    ��  �   T       �    ��  �   V       �    �  �   �       �    �\  �   U       �    4  �             ��  �   n           ��  �   }           �3  �   �           ��  �   �       "    ��  �   9       (    �% �          .    �  �   S       6    P8  �   j      ?    <�  �   k       J    Eh  �         �	    `" �           V    G�  �   W       ]    B~  �   H      h    ��  �   �       o    [�  �   �       v    ��  �   �       �    Bt  �          �    ڌ  �          �    (/  �   ]      �    Q�  �   X       �    �Y  �   �       �    v  �   �       �    >�  �   ]       �      �          �    �k  �   D      �    �- �          �    �^  �   �      �    6�  �   �       �    ��  �   �       B	       �           �    ��  �   9       	    )�  �   ;       	    ��  �   b       	    (% �          	    <"  �   �      	    A�  �   K       #	    n�  �   *       )	     �  �   K       0	    ��  �   �       8
    ��  �   /       8	    DU  �   r       @	       �           G	    0% �          '    ��  �   �       ?    j�  �   a       R	    7�  �         

    ��  �   S       [	    B  �   +       f    �W  �   �      i	    DS  �   �       q	    ��  �   l       �    �U  �         {	    ��  �   �       �	    ��  �   9       �	    �E  �   I       �	    ��  �   e      �	    `" �           �	    ��  �   9       �	    ��  �   K       !    ��  �         �	    v:  �         �	    ��  �   Z       �	    ԙ  �   6      �	    	�  �   9       �	    1�  �   �       �	    ��  �   2       [
    !�  �   �       �	    8% �          �	    �z  �   i      �	     �  �   �       �	    �R  �   �       �	    �  �   '      D
    ��  �   �       A	       �           
    @% �          	
    ��  �   S       
    �S  �   p       
      �   @      
    N   �           (
    ��  �   C      4
    d�  �   :       =
    ��  �   u      C
    ��  �   �       I
    ��  �   ]       P
    H% �          �     P �           Y
    0�  �   \      a
    C�  �   L       h
    U�  �   Y       �
       �           p
    ڍ  �   �       z
    Z�  �   7       
    P% �          �
    �  �   a       �
    d�  �   U       �    �@  �         �
    ��  �   �       R
    Q<  �   �      �
    H]  �   i       �
    ��  �   ;       �
    ݞ  �   3      �
    `   �   �      �
    �;  �   �       �
    
�  �   L       �
       �           �
    ��  �   U       �
    �A  �   9       �
    ^  �   �       �
    ��  �   '       �
       �           �
    �a  �   ^       E
    V�  �   �       
    ��  �   4           3�  �   a           ��  �   �           ��  �   9            ��  �   +      *    s�  �   =       0    ��  �   �      9    �  �   r       A    �\  �   U       M    ��  �   L       R    ��  �   O       lib/setup.asm HEADER_MAGIC HEADER_FLAGS header crt0.c launcher.c .LC60 .LC61 .LC62 .LC63 .LC64 .LC65 .LC66 .LC67 .LC68 wallpaper.c .LC0 .LC1 .LC2 .LC3 .LC4 .LC5 gui.c font8x16.c window.c bmp.c font.c border.c file.c cfs.c alloc_spin_lock pipe.c path.c memcmp.c memcpy.c memset.c strcasecmp.c strcat.c strchr.c strcmp.c strcpy.c strcspn.c string.c strlen.c strncasecmp.c strncmp.c strncpy.c strpbrk.c strrchr.c strsep.c strspn.c strtok.c last.1481 strstr.c strdup.c memmove.c strcoll.c strerror.c ctype.c tolower.c toupper.c stdio.c fopen.c fclose.c fflush.c fputc.c fgetc.c fgets.c fputs.c fread.c fwrite.c remove.c rewind.c fseek.c feof.c ftell.c vfprintf.c vf vsprintf.c vsnprintf.c sn_buf putchar.c sscanf.c perror.c vfscanf.c character _buf.1638 fvalue _buf.1650 ungetc.c getchar.c freopen.c tmpnam.c _tmpnam rename.c itoa.c i2hex.c malloc.c calloc.c free.c realloc.c lldiv.c strtol.c atoi.c atol.c strtoul.c exit.c getenv.c qsort.c qscmp qses qsexc qstexc qs1 system.c strtod.c ftoa.c _precision atof.c strtof.c strtold.c abs.c ltoa.c utoa.c srand.c errno.c gmtime.c localtime.c strftime.c clock.c math.c pow.c sqrt.c atan.c acos.c asin.c floor.c ceil.c exp.c locale.c signal.c setjmp.c _GLOBAL_OFFSET_TABLE_ longjmp read_directory_blk drawstring strcpy log sqrt setjmp clean_blk_enter put strtok_r stdout vsprintf ungetc pwd_ptr argv strerror utoa_r __m_i memmove __tm __realloc_r atol __window_puts getenv ceil errno floor strtold _infinity qsort fgets file_update file_read_block memcpy __window_clear BitMAP2 perror ltoa_r tolower system feof malloc remove fs_directory __window_putchar ldexp vsnprintf strtoul itoa __pipe__ stdgetc_r update_directory_entry _drawline fflush argc drawrect BitMAP eh_frame stdputc_r upath tell_r strncasecmp border write_r strtol user rename flush_r strrchr utoa calloc strtod rewind_r atof seek_r strcat read_directory_entry debug_o fseek __free_block_r open_dir ftoa stdin font8x16 __m_c _start obj_list __end strstr write_blk get_file_name atan2 signal strcoll strncmp write_sector draw_char_transparent pow strncpy put_pixel strcasecmp log10 _BLK_ realloc drawchar path_count open_file_r strtok remove_blk memcmp sscanf getfilename file_close pipe_write wp sigaction read_r file_write_block fread _ctype open_file addr search_blk_null strdup fopen sysgettmpnam localtime memset pwd main ftell srand fclose getchar close_r __data ptr_mouse2 __free_r update_window getkeyw _vsputs_r strcmp color remove_file __bss atan fgetc drawchar_trans strtof strcspn asin ltoa setlocale stderr create_file strsep getkey __malloc_r mouse fputc open_r A__ call_function getpathname strftime i2hex lldiv fwrite __window vfscanf rewind freopen pipe_read exit pipe_r __block_r atoi __heap_r assert_fn gmtime strspn ctr0 drawstring_trans strlen __code toupper wcl filename_cmp clock read_super_block abs strchr fputs acos strchrnul frexp vfprintf strpbrk read_sector free setpath  .symtab .strtab .shstrtab .text .data .got .got.plt .data.rel.local .bss .eh_frame .comment                                                                                  �           �                             !                �                                          '                �          h                              ,             h  �   h                                   5             �  �   �      �                              E             `" �   `"     �                             J              0 �    0                                    T      0                P     *                                                   0P     H*      
   �                 	                      xz     Z                                                   ҅     ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ELF          >       �   @       ��         @ 8  @                   �      �                                      �      �   �        @                   P      ` �    ` �    0       0             Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��  ���_ cole _          �      �            � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           I��H�D �   L�H��C �   H�H�   �   L�H�  �   L�#H�  �   L�+�   �����H��H��H��H��L�������UH��AWSH��@��H�����I�      L�H�}�H�u�H�U�H�M�L�E�L�M�H���������H�H�U�H�H��     H�E�H�H�E�H�`     H�H�`     H�H� H��H��     H�H��     H�H��H�P     H�H�`     H�H�@H��H�H     H�H�E�H�h     H�H�E�H�@     H�H�E�H��     H�H��     H�H��H�X     H�I�߸    H�e������H���H�p     H�    H���������H�H� H��H�x     H�H���������H�H� H��H���������H�H� H�։�I��H���������H��ЉE�E��I��H�ƻ������H��АH��@[A_]���UH��AWSH�� ��H�����I�%     L�H��     ��   H��     �   �    I��H���������H���H�E�H��jj h��� A�/ A�0  �  �    �   H���������H�<I��H�71������H���H�� H�E�H�E��@$H��     �)Љ�H�E��@(H��     �)Љ�H��     �4H��     �j�u�A���� A�    ��I��H��f������H���H��H�E�H�E�H��I��H��[������H���H�E�H��I��H��6������H���H�E�H��I��H�WU������H���H���������H�H� �   H���rH�E�H��H�v�������H�������UH��AWSH�� ��H�����I�{     L�H�}�H�E�H�ƿ    I��H��]������H��ЉE�}� t-�}�u(H���������H�<I�߸    H�ҟ������H������H�� [A_]���UH��AWSH����H�����I��     Lۉ}�H�u�H�E�� ��H�E��@9�sH�E��P#H�E��@9�r"H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@��u)H���������H�H��E�H�։�H� �������H���H�E�H�PH�E��@#��H�H�E�H�PH�E�H�@�U�H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  H�E��@��u0H���������H�H� H��t�E�����I��H��7������H��ЋE�H��[A_]���UH��H����H�����I��     L�H�}��E�    H�E�@��u]H�E�@'�PH�E�P'��H�E�P#H�E�@'9�r�H�E�H�PH�E�@'��H��H�H�E�H�PH�E�H�@� ���E��   H�E�@��tH�E�@��uiH�E�@#��u������ZH�E�P'H�E�@#9�r������AH�E�H�PH�E�@'��H�H�E�H�PH�E�H�@� ���E�H�E�@'�PH�E�P'�E�����UH��H����H�����I�|     L�H���������H�H� H�E��E�    H�E��@��uWH�E��P#H�E��@'9�w�    �AH�E�H�PH�E��@'��H�H�E�H�PH�E�H�@� ���E�H�E��@'�PH�E��P'�E�����UH��H����H�����I��     L�H���������H�H� H�E��E�    H�E��@��uXH�E��@'�PH�E��P'��H�E��P#H�E��@'9�r�H�E�H�PH�E��@'��H��H�H�E�H�PH�E�H�@� ���E��E�����UH��AWH��(��H�����I�)     L�H�}�H�u�H�U����u�    �(H�M�H�U�H��H��I��H���������H���H�E�H�E�H��(A_]���UH��AWSH�� ��H�����I��     L�H�}�H�}� u
������   H�}� tH�E؋@����tH�E��@"<t������zH�E؋@%�   ��u�    �cH�E؋@#H�U؋J�    ��E�H�E؋@��@��u�U�H�E؉�H��I��H��	������H���H�E�H��I��H��������H��ЉE�E�H�� [A_]���UH��AWSH����H�����I��     L�H�}�H�}� u������0H�E�H��H�9�������H���H�E�H��I��H�������H���H��[A_]���UH��AWSH�� ��H�����I�_     Lۉ}�H�u�H�}� u
�������  H�EЋ@��u
�    �  H�EЋ@��tH�EЋ@��tH�EЋ@��u!H�UЋE�H�։�H� �������H����y  H�EЋ@����unH�EЋP#H�EЋ�+  9�wYH�EЋ�+  ��tKH�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��E�U�H�EЉ�H��I��H�	������H����H�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U܈H�E�� ��H�EЋ@��9�r3H�EЋ@����H�EЉPH�E�f�   H�E�H��H�9�������H���H�EЋ@#�PH�EЉP#H�EЋP#H�EЋ�+  9�vH�EЋ�+  �PH�EЉ�+  H�EЋ@���H�EЉP�    H�� [A_]���UH��AWH��(��H�����I�D     L�H�}�H�}� u
������  H�E؋@��u
�    �v  H�E؋@��tH�E؋@��tH�E؋@��u"H�E�H��H�Z�������H��ЉE�E��0  H�E؋P#H�E؋�+  9�r
������  H�E؋@����ulH�E؋P#H�E؋�+  9�wWH�E؋�+  ��tIH�E؋@����H�E؉PH�E؋@#H�U؋r�    ���E�U�H�E؉�H��I��H�	������H���H�E؋@#H�U؋J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@� ���E�H�E�� ��H�E؋@��9�rH�E؋@����H�E؉PH�E�f�   H�E؋@#�PH�E؉P#�E�H��(A_]���UH��SH��H��H�����I�v     L�H�}ȉuĉU�H�M�H�}� u�    �y�E�    H�E�H�E��E�    �FH�E�H��H���������H��ЉE؃}��u�E�    �u��4H�E�H�PH�U��U؈�E��E��E��E��E�9�w��E�    �u�H��H[]���UH��SH��H��H�����I��     L�H�}ȉuĉU�H�M�H�}� u�    �l�E�    H�E�H�E��E�    �9H�E�H�PH�U�� ���E�H�U��E�H�։�H���������H��ЃE��E��E��E��E�9�w��E�    �u�H��H[]���UH��H����H�����I�     L�H�}�H�u��U�}�tZ�}�|�}� t�}�t�nH�E���H�E��P#H�E���H�E��P'�RH�E��@#H�U��H�E��P#H�E��@'H�U��H�E��P'�(H�E���+  H�U�)Љ�H�E��P#H�E��P#H�E��P'�H�E��@#H�U��J�    ��Љ�H�E�f��    ����UH��H����H�����I�$     L�H�}�H�}� u�    �	H�E��@#������UH��H����H�����I��     L�H�}�H�}� t7H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@����H�E��P������UH��H��(��H�����I�z     L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H��(��H�����I�%     L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H����H�����I��     L�H�}��E�_   �(�E�Hc�H�E�H�� < u�E�Hc�H�E�H��  �m��}� y����    ����UH��H����H�����I�g     L�H�}�H�E�H�E�H�E�H�E��H�E�� </uH�E�H��H�E�H�E�H�E�� ��u�H�E�����UH��H��0  ��H�����I��     L�H������H������H������H�E�H������H�E�H������H�E��E�    �?H�E�� ��u�E�Hc�H�E�H��  �H�E�H�PH�U��U�Hc�H�U�H�� ��E��}�_~��E�    �-H�E�H�PH�U��H�E�H�PH�U�� 8�t�   ��E��}�_~͸    ����UH��SH�� ��H�����I�     L�H�}�H�u�H�E؋PH�E؋@ЉE�E�H�U����H��     H�H�¾   H�z�������H��ЉE�}� t
�������   �E�    ��   �E�%�  ��H��     ��H؋���uf�E�%�  ��H��     ��H��������E�H�U����H��     H�H�¾   H���������H��ЉE�}� t������r�E��m�E�%�  =�  uE�E��E�H�U����H��     H�H�¾   H�z�������H��ЉE�}� t�������E�H�E؋@$9E����������H�� []���UH��H����H�����I��     L؉}��u�H�U�H�M�    ����UH��AWSH��0��H�����I�S     Lۉ}�H�u�H�U�H�EȋPH�Eȋ@ЉE�H�Eȋ@ �E܉E�ЉE�   �    H��     H�<I��H�q������H����E�    �B�U�E�Љ�H�EЋ ��H��     H��   H���������H��ЉE��}� u�E�H�EȋP �E�9�w���H��0[A_]���UH��H����H�����I�m
     L�H�}�H�u�H�U��R��H�U����H�U�H��H��   I�z�������J� ������UH��AWSH��`��H�����I�
     L�H�}�H�u�H�U�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�E�H�E�H�E�H��I��H�'������H��ЉE�H�E��@,�E��9  H�E�H�E��H�E�� </uH�E��  H�E��H�E�H�E�� ��u׋U�H�E��@ H�M��	��H�M���H�z�������H��ЉE؃}� t#H�E�H��I��H�#�������H��и    ��   �E�    �f�E���Hc�H�E�H�H�E�H�E��@a��t5H�E��@b����@��t#H�E�H�U�H��H��H���������H��ЉE���E������}� t�E��}�?~����}� u+�}�?%H�EЋ@k�E�H�E��@ �E؉E�ЉE�m��	�E�    �
�}� �����H�E�H��I��H�#�������H��ЋE�H��`[A_]���UH��AWSH��P��H�����I��     L�H�}�H�u�H�U��M�L�E�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�Eغ    �    H��I��H�q������H��ЋU�H�E��@ H�M��	��H�M؉�H�z�������H��ЉE�}� t#H�E�H��I��H�#�������H��и������   �E�    �T�E���Hc�H�E�H�H�E�H�E��@a��t#H�E�H�U�H��H��H���������H��ЉE���E������}� t�E��}�?~����}� u:�}�?4�E���Hc�H�E�H�H�EȺ�   H��H��I��H��p������H�����E�����H�E�H��I��H�#�������H��ЋE�H��P[A_]���UH��AWSH��P��H�����I�-     L�H�}�H�u�H�U�H�E���C  ��u
������	  H�E���C  ��@v/H��������H�<I�߸    H�ҟ������H��Ҹ������  H�E��PH�E��@ЉE�H�E���?  H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�Eغ    �    H��I��H�q������H��ЋU�H�E��@ H�M��	��H�M؉�H�z�������H��ЉEԃ}� t!H�E�H��I��H�#�������H��ЋE��  H�E���C  ��H��H��H�E�H�H�E�H�EȺ`   �    H��I��H�q������H���H�E�H��+H��H���������H���H��H�E�H��H��I��H��s������H����E�    �"H�UȋE�H����uH�UȋE�H�� �E��}�_~�H�E��@` H�E���+  H�EȉPo�U�H�E��@ H�M��	��H�M؉�H���������H��ЉE�H�E�H��I��H�#�������H��ЋE�H��P[A_]���UH��AWSH��`��H�����I��     L�H�}�H�u�H�U��S  I��H���������H���H�E�H�EкS  �    H��I��H�q������H���H�E��PH�E��@ ��H�EЉP�    I��H���������H���H�U�H�BH�E��PoH�EЉ�+  H�E��PH�EЉ�/  H�E��P H�EЉ�3  H�E��H�EЉ�G  �    I��H���������H���H�U�H��K  H�E�H��K  �    �    H��I��H�q������H���H�E��@k�E�    I��H���������H���H�E��E������E�    �E�    ��  �   I��H���������H���H�U�H��K  �M�Hc�H��H�H�H�E�H��K  �U�Hc�H��H�H� H�E�H�E��   �    H��I��H�q������H����E�    �<  H�E��@ �E��H�E��@�H�E��P�E�H�H�4�    H�E�H�ʉH�EЋ�;  �PH�EЉ�;  �E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E�;E�ts�E�H�U����H�U�H��H�¾   H�z�������H��ЉE��}� t:H�E�H��I��H�#�������H���H�E�H��H�������H��и    �   �E��E�H�E��@�����E�    ��U�E�H��    H�E�HЋ �E�}��u	�E�������E��}��  ������}��t�E��}��  � �����H�E�H��I��H�#�������H���H�E�H��`[A_]���UH��AWSH��p  ��H�����I�N      L�H������H�������   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H������H�E�H��H��I��H��$������H���H�U�H�E�H��H��I��H��'������H��п�   I��H���������H���H��     H�H��     H���   �    H��I��H�q������H��п   I��H���������H���H�E�H�EȺ   �    H��I��H�q������H���H�E�H�E�H�E��   �    H��I��H�q������H����E�    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ ���    Hǅ���    Hǅ���    Hǅ���    Hǅ ���    Hǅ(���    Hǅ0���    Hǅ8���    Hǅ@���    HǅH���    HǅP���    HǅX���    Hǅ`���    Hǅh���    Hǅp���    Hǅx���    H�E�    H�E�    H������H������H��H��I��H��s������H���������<wt������<au�E�   H�E��@   H�E��     H�U�H�E�H��H��H���������H��ЉE�}� t_H��     H�H��I��H�#�������H���H�E�H��I��H�#�������H���H�E�H��I��H�#�������H��и    �  H�E�H�U�H�M�H�E�H��H��H���������H��ЉE��}� u_H��     H�H��I��H�#�������H���H�E�H��I��H�#�������H���H�E�H��I��H�#�������H��и    �  H�EȋU��P,H��     H�H�M�H�U�H�u�I�ȹ    H��H���������H��ЉE�}����   �}� tqH��     H�H������H�U�H�u�A�    H��H��������H���H��     H�H������H�U�H�u�I�ȹ    H��H���������H��ЉE�}� ��   H��     H�H��I��H�#�������H���H�E�H��I��H�#�������H���H�E�H��I��H�#�������H��и    ��  �}� t_H�E�H��I��H�#�������H���H��     H�H��I��H�#�������H���H�E�H��I��H�#�������H��и    �r  H��     H�H�U�H�M�H��H��H�!�������H���H�E�H�}� ��   H��     H�H��H�E�H��+�`   H��H��I��H��p������H���H�E�H��+H��H�$�������H���������<wt������<+t������<au
H�E��@"�H�E��@"H�E��@   H�EȋP,H�E���?  H��     H��PsH�E���C  ������<auH��     H��PoH�E��P#H�E�H��I��H�#�������H���H��     H�H��I��H�#�������H���H�E�H��I��H�#�������H���H�E�H��p  [A_]���UH��AWSH��@��H�����I��      L�H�}��   I��H���������H���H�E�H�E�   �    H��I��H�q������H���H�E�H�E�H�E�   �    H��I��H�q������H���H�E��@   H�E��     H�U�H�E�H��H��H���������H��ЉE܃}� t H�E�H��I��H�#�������H��и�����AH�U�H�M�H�E�H��H��H���������H��ЉE�H�E�H��I��H�#�������H��ЋE�H��@[A_]���UH��AWSH�� ��H�����I���      L�H�}�H�E�H�@H��I��H�#�������H����E�    �TH�E�H��K  �U�Hc�H��H�H� H��t?H�E�H��K  �U�Hc�H��H�H� H��I��H�#�������H��ЃE��}��  ~���H�E�H��K  H��I��H�#�������H���H�E�H��I��H�#�������H���H�E�    �    H�� [A_]���UH��H�� ��L�����I���      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H�z�������I� ������UH��H�� ��L�����I��      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H���������I� ������UH��AWSH��   ��H�����I�(�      L�H��x���H��p�����l����   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H��x���H�E�H��H��I��H��$������H���H�U�H�E�H��H��I��H��'������H��п   I��H���������H���H�E�H�EȺ   �    H��I��H�q������H���H�E�H�E�H�E��   �    H��I��H�q������H���H�E��@   H�E��     H�U�H�E�H��H��H���������H��ЉE��}� t_H��     H�H��I��H�#�������H���H�E�H��I��H�#�������H���H�E�H��I��H�#�������H��и�����-  H�E�H�U�H�M�H�E�H��H��H���������H��ЉE��}� u_H��     H�H��I��H�#�������H���H�E�H��I��H�#�������H���H�E�H��I��H�#�������H��и�����  H�EȋU��P,H�EȋPH�Eȋ@ЉE�H�EȋP,H�Eȋ@ �ЋE�ЉE��    I��H���������H���H�E�H�E��    �    H��I��H�q������H��ЋU�H�Eȋ@ H�M��	��H�M���H�z�������H��ЉE��E�    �E�    �   �E���Hc�H�E�H�H�E��E�;�l���}~H�E��@a��ta�E���Hc�H��p���H�H�E���   H��H��I��H��p������H��ЋE���Hc�H��p���H�H��H�$�������H��ЃE����E��}�?�e�����H�E�H��I��H�#�������H���H�E�H��I��H�#�������H���H�E�H��I��H�#�������H��ЋE�H�Đ   [A_]���UH��AWSH��`��H�����I�<�      L�H�}�H�u�H�U�H�M�D�E�H�E�H�E�H�Eغ�   �    H��I��H�q������H���H�E�H��H���������H���H��H�E�H��H��I��H��s������H����E�    �"H�U؋E�H����uH�U؋E�H�� �E��}�_~�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉEп    I��H���������H���H�E�H�EȺ    �    H��I��H�q������H��ЋU�H�E��@ H�M��	��H�Mȉ�H�z�������H��ЉEă}� t!H�E�H��I��H�#�������H��ЋE���  �E�    �$�E���Hc�H�E�H�H�E�H�E��@a��t�E��}�?~���H�E��@a���G  �}�?�=  �U�H�E؉PsH�E��@a��E���H�E؈PbH�U�H�E�H��H��H���������H���H�U؉BkH�E؋@k���uOH�E�H��H�$�������H�<I�߸    H�ҟ������H���H�E�H��I��H�#�������H��и   ��   �E���@��t$H�E؋@kH�U�H�M�H�Ή�H���������H���H�M�H�E຀   H��H��I��H��p������H��ЋU�H�E��@ H�M��	��H�Mȉ�H���������H��ЉEĐH�E�H��I��H�#�������H��и    �JH�E�H��I��H�#�������H���H�E�H��H�H�������H�<I�߸    H�ҟ������H��Ҹ����H��`[A_]���UH��AWSH��P��H�����I���      Lۉ}�H�u�H�U��    I��H���������H���H�E��E�    �E��E��E������E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E��E܋E�;E���   �}� tV�E�H�U����H�U�H��H�¾   H���������H��ЉẼ}� t#H�E�H��I��H�#�������H��и�����?  �E�H�U����H�U�H��H�¾   H�z�������H��ЉẼ}� t#H�E�H��I��H�#�������H��и������   �E��E�E��E��E�   H�E��@�����E�    ��U�E�EȋE�H��    H�E�HЋ �E�E�H��    H�E�H��     �}��uL�E�H�U����H�U�H��H�¾   H���������H��ЉE̐H�E�H��I��H�#�������H��ЋE��6�E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��Y���H��P[A_]���UH��AWSH��   ��H�����I���      L�H��h����   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H��h���H�E�H��H��I��H��$������H���H�U�H�E�H��H��I��H��'������H��п   I��H���������H���H�E�H�E��   �    H��I��H�q������H���H��p���H�E�H�E��   �    H��I��H�q������H���H�E��@   H�E��     H�U�H�E�H��H��H���������H��ЉE�}� t<H�E�H��I��H�#�������H���H�E�H��I��H�#�������H��и    ��  H�E�H�U�H�M�H�E�H��H��H���������H��ЉE��}� u<H�E�H��I��H�#�������H���H�E�H��I��H�#�������H��и�����d  H�E��U��P,H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE��    I��H���������H���H�E�H�E��    �    H��I��H�q������H��ЋU�H�E��@ H�M��	��H�M���H�z�������H��ЉE�}� tSH�E�H��I��H�#�������H���H�E�H��I��H�#�������H���H�E�H��I��H�#�������H��ЋE��l  �E�    �   �E������E���Hc�H�E�H�H�E�H�E��@a��t!H�E�H�U�H��H��H���������H��ЉE�}� u9H�E��@a �U�H�E��@ H�M��	��H�M���H���������H��ЉE�}� ��E��}�?�k����}� tPH�E�H��I��H�#�������H���H�E�H��I��H�#�������H���H�E�H��I��H�#�������H��ЋE��uH�E��@kH�U�H�M�H�Ή�H�������H��ЉE�H�E�H��I��H�#�������H���H�E�H��I��H�#�������H���H�E�H��I��H�#�������H��ЋE�H�Đ   [A_]���UH��H����H�5����I�)�      Lމ}�E�E��}� u�E��   �E����rH��     H�H��     H�����UH��H����H�����I���      L�H�}��   H�E�H���r�����UH��AWH����H�����I���      L�H��     H�H�U�H��     H�    H�P       �    H�M�   �    H��I��H�q������H��ѐH��A_]���UH��AWSH��P��H�����I��      Lۉ}��u��}� u
�    ��  H��     H�H=�   v%H���������H�<I�߸    H�ҟ������H��ҐH�P       ���u�H�P       ��PH�P       ��E����E�E�%�  ��t�E��E�    �E�    �E�    �}� t�E��   �E�   �K  �}��  �=  H��     H�H�E�H�E�    �E�    �  H�E؋@����   H�E؋@9E���   H�E�H�H�E؋@��H�H�E�H�E؋@+E���H�E؉PH�E؋P�E��H�E؉PH�E�H�E�H��     H�H�E��E�    �mH�E؋@��tH�E��E��WH�E�H�E�H�E�H�E�H�E�H�@H�PH�E�H�PH�E��@   H�E�H�U�H�H�E��U��PH�E�H�U�H�P�E���!�}��   ~��H�E��E��}��   ������E�   ���}� ��   H��     H�H�E��E�    �~H�E؋@��tH�E��E��hH�E�H�E��E��H��������H���H�E�H�E�H�U�H��E��E���H�E��PH�E��U��P�E���+E���H�E��PH�E�H�@   ��}��   �u���H�P       �    H��     H�H�PH��     H�H�E�H��P[A_]���UH��SH��(��H�����I���      L�H�}�H�}� ��  �H�P       ���u�H�P       ��PH�P       �H�E�H�E�H��     H�H�E��E�    �M  H�E�H� H9E�tH�E��E��2  H�E�H�E�H��     H�H�P�H��     H�H�E؋@��uH�E�H��H�,������H����   H�E؋@��uH�E�H�@H�E�H�E�H�@H�P�H�E�H�PH�E�H�@H��tH�E؋@����   H�E�H�@H��uRH�E�H� H��H�,������H���H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    ��}��   �������H�P       �    ��H��([]���UH��AWH��H��L�����I���      M�H�}��u�H�E�    �E�    H�}� u�E��   ��H��������I� ���8  �H�P       A� ��u�H�P       A� �PH�P       A� H��     I� H�E�H�E�H�E��E�    �   H�E�H� H9E�t
H�E��   H�E�H�E��E�   H�E��P�E��=   v@H��     I� �U�H�E�H��H���������I�< M�Ǹ    I�ҟ������M�A����H�E�H� H�E�H�E��P�E��H�E��P�E��}��   �X���H�P       A�     �}� u�E��   ��H��������I� ���H�E�H��HA_]���UH��H�� ��H�����I�>�      L�H�}�H�u��E�    H�E�H�E��   H�E�� ��H�E��@9�sH�E��P#H�E��@9�rH�E��@#    H�E�f�   H�E�H�PH�E��@#��H�H�E�H�PH�E�H�PH�U�H�U�H�R� �H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  �E��}��E����E�����UH��H�� ��H�����I�>�      L�H�}�H�u��E�    H�E�H�E�H�E��@'�PH�E��P'H�E��P'H�E��@9�rH�E��@'   �H�E��P#H�E��@'9�r�H�E��@'�P�H�E��P'�JH�E�H�PH�E��@'��H�H�E�H�PH�E�H�PH�E�H�HH�M���H�E��@'�PH�E��P'�E��}�~��E�����UH��AWSH��0��H�����I�W�      L�H�}�H���������H�H� H�E�H�E�H�E�H�E�H��I��H�vv������H��ЉE�H�E�H��I��H�vv������H��ЉE؋U܋E��=   ~
������   H�E�� </uH�E��E�H�HE�H�m�H�E�� </tH�E�H�E�H�PH�U�� /�H�E�H�U�H�E�H��H��I��H��s������H���H�E�H��I��H�vv������H��Љ�HE�H�m�H�E�� </u	H�E��  �H�E�H�E��  �    H��0[A_]���UH��AWSH����H�����I��      L�H���������H�H� H��I��H�vv������H��Ѓ�w
�    �   H���������H�H� H�E�H�E�H��I��H�vv������H��Љ�HE��H�E�H�P�H�U��  H�E�� </u�H���������H�H� H��I��H�vv������H��Ѓ�vH�E��  �    H��[A_]���UH��AWSH��0��H�����I��      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
�    ��  H�E�H��I��H�vv������H��ЉE�E�H�H�P�H�E�H�� </u�E�H�H�P�H�E�H��  �}� 
�    �  �}���   H�E�H��� <:u%H�U�H�E�H��H��I��H��s������H����K  H��������H�<I��H���������H���H��H�E�H��H��I��H��s������H���H�E�H��I��H�vv������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H��s������H����   H��������H�<I��H���������H���H��H�E�H��H��I��H��s������H���H�E�H��I��H�vv������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H��s������H���H�E�H��0[A_]���UH��H����H�����I���      L�H�}�H�E�H�E�H�}� u�    �+�E�    �H�E�� </u�E�H�E�H�E�� ��u�E�����UH��AWSH��0��H�����I�n�      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
������   H�E�H��I��H�vv������H��ЉE�E�H�HE�H�m��H�E�� </tH�m�H�E�� ��t�E�P��U�����H�E�H�U�H�E�H��H��I��H��s������H���H�E��  �    H��0[A_]���UH��H��0��H�����I���      L�H�}�H�u��U܉M�L�E�H���������H�H� H�E��E�H9E�}?H�E��@��H9E�}0H�E�H�E��E�H�E�H��H�E�H�H��    H�E�HE؉������UH��SH��@��H�����I���      Lۉ}ԉuЉỦM�L�E�L�M�f�E�  H�E�H�@H�E�H�E��@�E�}�u�E�    �E�    �   f�E� H�E��@�EȉE��H�H� H�E�H�� f�E�H�E�� ���E��J�E�f#E�f��t5�UЋE��Hc��UԋE��H�H�}��M�U�I��H��H�k(������H���f�e�m��}� y��E�H�E��@9E��b�����H��@[]���UH��AWSH��0��H�����I���      Lۉ}܉u؉UԉM�D�E�L�M��E�    �X�E�    �CH�E�L��   �M�H�E��P�u؋E��Hc��}܋E��H�H��I��H�k(������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I�,�      Lۉ}܉u؉UԉM�D�E�L�M��E�    �p�E�    �[H�E�H��   �E��E�i��E��A��H�E��P�M؋E��Hc��M܋E��H�I��D��H��I��H�k(������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I�e�      Lۉ}܉u؉UԉM�D�E�L�M��}� �[  �}� �Q  �E�    �>H�E�L��   �M�H�E��P�E�Hc��}܋E��H�H��I��H�k(������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E����Hc��}܋E��H�H��I��H�k(������H��ЃE��E�;E�|��E�    �AH�E�H��   �M�H�E��P�u؋E��Hc��E�H�I��H��I��H�k(������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E��Hc��}܋E����H�H��I��H�k(������H��ЃE��E�;E�|���H��0[A_]���UH��AWSH��@��H�����I���      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}��  �E�    ��   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��   �E�f#E�f��tDH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�k(������H����BH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�k(������H���f�e�m��}� �[����E�H�E��@9E��	�����H��@[A_]���UH��SH��8��H�����I�S�      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H�6-������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I���      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}���   �E�    �   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��W�E�f#E�f��tBH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�k(������H���f�e�m��}� y��E�H�E��@9E��T�����H��@[A_]���UH��SH��8��H�����I�x�      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H�\/������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I���      L�H�}ȉuĉU��M�D�E�D�M�H���������H�H� H�E�H�E�H   � �? �    H��I��H�q������H����E�    �U�H�E��P4�UH�E��P8�UH�E��P<H�E��@H   H�E��@L   H�E��P<H�E��PP�UH�E��PTH���������H�H��H�E�H�PXH�E��@D    H�E��PDH�E��P@�U�H�E��P�U�H�E��P�U�H�E��P �U�H�E��P�U H�E��P`�} u�E�   H�E��@�P�H�E��P(H�E��P�E�)ЍP�H�E��P$H�E��@0   �E����H�E��P,H�E��@��H�E��@��H�E�I���Ѻ    �    I��H��A������H���H�E��@4��H�E��@����H�E�I��A�ȹ   �   �   H�*������H��Ѓ}� u:H�E��@����H�E�I��A���� �   �   �   H�*������H����8H�E��@����H�E�I��A���� �   �   �   H�*������H��Ѓ}� t}H�E��@����H�U��E�I��A���� ����   �   H�*������H���H�E��@4��H�E��@���ƋE��H�U�I��A�ȹ   ��ƿ   H�*������H���H�E��@8A��H�E��@$��H�E��@(��H�E��@,��H�E��@0��H�E�I��H�*������H���H�E�H��I��H�vv������H������E�H�E�H�pHH�E��@��E܉������)Љ�H�E�H���u�I��A���� ������   ��H��H�{0������H���H��H�E��@����H�E�I��A�    �   �   �   H��+������H���H�E�H�PHH�E��@��H���u�I��A���� ������   �ƿX   H�\/������H���H��H�E�H�PHH�E��@��(H���u�I��A���� ������   �ƿ-   H�\/������H���H��H�E�H�e�[A_]���UH��AWSH��0��H�����I�6�      L�H�}�H�u�H�E��P0H�E��@Ѓ�P�E�H�E��P,H�E��@Ѓ��E��E�P   �E�   �E�    �E���� H�E�H��I��H�vv������H��ЉE�H�E�L�@H�M؋U܋E���������p��E�<�E��������ƋE���)ƋE��H�E�H���u�M��A�ȉщ�H��H��.������H���H���H�e�[A_]���UH��H����H�����I�2�      L�H�}��   H�E�H���r�����UH��H����H�����I���      L�H�}������UH��H����H�����I���      L�H�}�H�U��BD    H�U��JDH�U��J@H�U��R8A��H�U��R$��H�U��R(A��H�U��R,��H�U��R0��H�U�I��D��I�*������J��А����UH��SH��(��L�����I�@�      Mډ�f�E�H���������I�H� H�E�H���������I�H��H�E�H�PXH�E�@(�P�H�E�@H���к    ��E�H�E�@$�P�H�E�@L���к    ��E�H�E�P<H�E�PPH�E�PD�E�9�rH�E��@D    H�E�@@�PH�E�P@H�E�P@�E�9�r9H�E��@D    H�E�PDH�E�P@H�E�H��H�&7������I����E��  f�}���   H�E�@D����   H�E�@D�P�H�E�PDH�E�H�xHH�E�pTH�E�@PH�U�J,H�U�RLA��H�U�R@A��ʃ���H�U�J0H�U�RHA��H�U�RDA��ʃ�A��H���u�I��A������D�޿    H�6-������I���H����   f�}�	uH�E�@D�PH�E�PD��   f�}�
u!H�E��@D    H�E�@@�PH�E�P@�   f�}���   H�E�H�xHH�E�pTH�E�PPH�E�H,H�E�@LA��H�E�@@A��ȃ���H�E�H0H�E�@HA��H�E�@DA��ȃ�A���E�H���u�I��A���щ�D�މ�H�6-������I���H��H�E�@D�PH�E�PD�E�H�]�����UH��H����H�����I�{�      L؉}�H���������H�H� H�E��U�H�E��P<�����UH��SH��(��H�����I�1�      L�H�}�H�}� t=H�E�H�E��&H�E�H�PH�U�� f�����H��7������H���H�E�� ��u���H��([]���UH��AWSH��P��H�����I���      L�H�}��u��U��M�L�E�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H��������H�<I�߸    H�ҟ������H��Ҹ�����6  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H��������H�<I�߸    H�ҟ������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�.�������H�<I�߸    H�ҟ������H��Ҹ   ��   �E�    �   �E�    �   �}� tNH�E�H��   H�E��P�M��E���E��Hc��M��E���E��H��M�I��H��I��H�k(������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�k(������H��ЃE��}� �U����E��}� �;����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��P��H�����I���      L�H�}��u��U��M�D�E�L�M�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H��������H�<I�߸    H�ҟ������H��Ҹ�����3  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H��������H�<I�߸    H�ҟ������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�.�������H�<I�߸    H�ҟ������H��Ҹ   ��   �E�    �   �E�    �   �}� tKH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�k(������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�k(������H��ЃE��}� �X����E��}� �>����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��0��H�����I���      Lۉ}܉u؉U�H�M��E�    �   �E�    �t�U�������E��H���������H�Hڋ��E�}� tBH�E�H��   H�EȋP�MԋE��Hc��M؋E��H��M�I��H��I��H�k(������H��ЃE��}�~��E��}��o�����H��0[A_]���UH��AWSH��@��H�����I��      Lۉ}̉uȉUĉM�L�E��E���� �E�``` �E���� �EĉE��ẺE܋E��E؋EȉEԋE؍P��E��xH�M��E�I��A�    �   ��I��H��+������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H��+������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H��+������H��ЋEԍP��E܍pH�M��E�I��A�    �Ѻ   ��I��H��+������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H��+������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H��+������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H��+������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H��+������H��ЋEԍP��E܍p�M��E�ȃ�H�M�I��A�    �Ѻ   ��I��H��+������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H��+������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H��+������H��ЋE؍P��M܋E�ȍp��E���H�M�I��A�    �   ��I��H��+������H��АH��@[A_]���UH��AWSH��0��H�����I��      Lۉ}܉u؉UԉM�D�E�D�M�H�} u
�    ��  �H   I��H���������H���H�E�H�}� u
�    ��  H�E�H   �    H��I��H�q������H���H�UH�E�H�P@H�E�U�PH�E�P0�E��H�E�PH�E�P,�E��H�E�PH�E��    H�E�P(�E�9�wH�E�P(H�E�P�
�U�H�E�PH�E�P$�E�9�wH�E�P$H�E�P�
�U�H�E�P�U�H�E�P�U�H�E�P H�E��@0    H�E�@0��I��H���������H���H��H�E�H�P8H�E�H�@8H��t.H�E�@0H�U�H�R8H�щ¾    H��I��H�q������H���H�E�@ ��H�E�@��H�E�@��H�E�@��H�E�@L�MA����I��H�*������H���H�E�@��H�E�@��H�E�@��H�E�@L�MA�������I��H��+������H���H�E�H��0[A_]���UH��AWSH�� ��H�����I���      L�H�}�H�E�H�@@H�E�H�E؋@ A��H�E؋@��H�E؋@��H�E؋@��H�E؋@��H�E�I��I��H�*������H���H�E�H��H��J������H��АH�� [A_]���UH��AWSH�� ��H�����I��      L�H�}�H�}� u
������z  I�߸    H�x�������H��҉E�}���   I�߸    H�x�������H��҉E�}�[��   I�߸    H�x�������H��҉E�}�Ct�}�Dt'�GH�E؋P,H�E؋@49�s1H�E؋@,�PH�E؉P,�H�E؋@,��tH�E؋@,�P�H�E؉P,����H�E�H��H��J������H��и    �  H�E�H�P8H�E؋@,��H�H�E��}� �C  H�E؋P,H�E؋@09��-  H�E��@    �}���   H�E؋@4��tkH�E؋@,��t`H�m�H�E؋P4H�E؋@,)�H�E�H�HH�E�H��H��I��H�B~������H���H�E؋@,�P�H�E؉P,H�E؋@4�P�H�E؉P4�   H�E��@   �~H�E؋P,H�E؋@49�t4H�E؋P4H�E؋@,)�H�E�H�HH�E�H��H��I��H�B~������H��ЋE��H�E��H�E؋@,�PH�E؉P,H�E؋@4�PH�E؉P4H�E��@   H�E�H��H��J������H���H�E؋@����u*H�E�H��H��J������H���H�E؋@����H�E؉P�    H�� [A_]���UH��AWSH��@��H�����I�E�      L�H�}�H�E�H�@@H�E�H�E�H�@8H�E��E�    f�E�  H�E��@��uH�E��@    �  �E�    �  �E�    �E�    ��   �}� ueH�E��P4�E�9�vH�E�H�PH�U�� f�f�E��f�E�  f�}�
uf�E�  �E�   H�E��P,�E�9�u�U�H�E��P$�U�H�E��P(�E�f�}� teH�E�H�xHH�E��p H�E��PH�E��H�E��A��H�E��H�E��A���E�H���u�I��A����D��D�։�I��H�6-������H���H���E�H�E��P�E�9������E�H�E��P�E�9������H�E�H�xHH�E��p H�E��@H�U��JH�U��R(�A��H�U��JH�U��R$�A��H���u�I��A����D��D�ֿ_   I��H�\/������H���H��H�e�[A_]���UH��AWSH��@��H�����I�B�      L�H�}�H�E��@ �E�H�E��@�E�H�E��@�E�H�E��@�E�H���������H�H� � �E�H���������H�H� �@�E�H���������H�H� �@�E̋EЃ����X  �E�;E�~Q�E���9E�~F�U�E��9E�}9�E��P�E��9E�})�E�+E��E�+E�։�I��H� W������H�����   �E�;E���   �E�;E���   �U�E��9E���   �U��E��9E���   H���������H�H� � ��H�E��@ )ЉE�H���������H�H� �@��H�E��@)ЉE��aH���������H�H� � +EȉE�H���������H�H� �@+EĉE�}� y�E�    �}� y�E�    �U�H�E��P �U�H�E��PH���������H�H� �@����u�I�߸    H�
V������H��ҐH��@[A_]���UH��AWSH��@��H�����I�$�      L�H�}�H�u�H�UȉM�D�E�D�M��P  I��H���������H���H�E�H�E�P  �    H��I��H�q������H���H�E�H��I��H�vv������H��ЉE�}�~�E�   �U�H�E�H�H0H�E�H��H��I��H��p������H���H�E��    H�E��U�P�U�H�E��P�E�����H�E��P�U�H�E��P�UH�E��PH�U�H�E�H�P(H�E�H�PHH�E��@����H�E��@����H�E�H��0H���u�I��A���� �    ��H��I��H��.������H���H��H�E�H�U�H��H�e�[A_]���UH��AWSH��0��H�����I���      L�H�}�H�uЉU�H�E؋@$��H��H��H�H��H�PPH�E�H�H��H�E�H�E؋@$�HH�U؉J$H�U؉�H��H��H�H��H�H�PP�ẺH�E�H��I��H�vv������H��ЉE�}�~�E�   �U�H�M�H�E�H��H��I��H��p������H��и    H��0[A_]���UH��AWSH��P��H�����I���      L�H�}��E�    �E�����H�E�H�@(H�E�H�E�H�PHH�E��@����H�E��@����H�E�H��0H���u�I��A���� �  � ��H��I��H��.������H���H��H�E�H�PHH�E��@����H�E��@��H���u�I��A���� �  � ���H�H�������H�<I��H�{0������H���H��H�E؋P0H�E��@ЉE�H�E؋@,�E��E�d   �E�   �EĀ�� �E�    �H���������H�H� �@����u�H�E��@$���A  H�E��P$�E���A��H�}؋MċŰuЋE�I��A��D�щ�I��H�*������H����E�    �  H���������H�H� � ��H�E؋@ )ЉE�H���������H�H� �@��H�E؋@)ЉE�H���������H�H� �@�E�E�Hc�H��H��H�H��H�PPH�E�H�H��H�E��E�;E���   �E��E��E�Ѓ�9E���   �UԋE��9E�}�E��E��E�E��9E�}gH�E�H�xH�MċE��E��E�ЍP�EԍpH�E�H���u�I��A�ȹ����H��I��H��.������H���H���E��E�m��E����tZ�nH�E�H�xH�MċE��E��E�ЍP�EԍpH�E�H���u�I��A�ȹ    H��I��H��.������H���H���E������E�H�E��P$�E�9��[����E�����A����}��t5H�M��E�Hc�H��H��H�H��H�H��P� ��I��H�A^������H����E�   �H���������H�H� �@����u�H�E�H�PHH�E��@����H�E��@����H�E�H��0H���u�I��A���� �    ��H��I��H��.������H���H���E�H�e�[A_]���UH��AWSH����H�����I���      L�H�}�H�X       H�    H�`       H�    I�߸    H��_������H���H�h       �    H�}� t'H�E� ��H�h       �H�`       H�E�H��    H��[A_]���UH��AWH����H�����I��      L�H�h       �����   ����   ��t
��tA�   H�`       H�H����   H�`       H�H��I��H��G������H����yH�`       H�H��tbH�M�������H�<I�׸    H�ҟ������H����?H�`       H�H��t+H�`       H�H��I��H�i������H����������    H��A_]���UH��AWSH��@��H�����I�Ѩ      Lۉ}��u�H���������H�H� H��t�}� x�}� y&�H���������H�H� �@����u������#  H�E�    H�E�    �E�    �E�    �E�    �E�    �   H��     �E�H�H�H��H�E�H�E�H��� �E�H�E�H��� �E�H�E�H��� �E�H�E�H��� �EċEԉE܋E�;E�~"�E�;E�~�UЋE��9E�}�ŰE��9E�|&�E��E�Hc�H���������H�H� H9��^������E�Hc�H���������H�H� H9�u&�H���������H�H� �@����u������  H�E� ���V  ����  ����  ���n  ��t����   �[  H��     �E�H�H�H��H��H�X       H�H�X       H�H�@(H�E�H�X       H��@��I��H�A^������H���H�X       H�H��I��H�:Q������H��ЉE���  H��     �E�H�H�H��H��H�`       H�H�`       H�H�@@H�E�H�`       H��@��I��H�A^������H����E�    H�h       �   �H���������H�H� �@����u��]  H��     �E�H�H�H��H��H�`       H�H�`       H�H�@@H�E�H�`       H��@��I��H�A^������H����E�    H�h       �   �H���������H�H� �@����u���   H��     �E�H�H�H��H��H�`       H�H�`       H�H�@@H�E�H�`       H��@��I��H�A^������H����E�    H�h       �   �H���������H�H� �@����u��*�H���������H�H� �@����u��E�    ������I�}� t>��H�E�� ��u�H�E�� �PH�E��H�E�H��H��\������H���H�E��     �    H��@[A_]���UH��AWSH����H�����I�0�      L�H�}�H���������H�H� H��u*�   �    H��     H�<I��H�q������H���H���������H�H� H=�   ~�    �LH���������H�H� H�HH���������H�H�
H�U�H��     H�H��H���������H�H� H��[A_]���UH��AWSH�� ��H�����I�P�      L�H�}�H�E�    H�E؋@8A��H�E؋@$��H�E؋@(��H�E؋@,��H�E؋@0��H�E�I��I��H�*������H����E�    �   H��     �E�H�H�H��H�E�H�E�� ��tWH�E�� ��uOH��     �E�H�H�H��H��H�`       H�H�`       H�H��I��H�NG������H��������E��E�Hc�H���������H�H� H9��\�����H�� [A_]���UH��AWSH�� ��H�����I��      Lۉ}�H�u�H�E�H��I��H��L������H��и    H�_������H��҉E�E�H�� [A_]���UH��H����H�����I���      L؉}�H��     ���	v5H��     �D    H��     �    H��     �D    H��     ��JH��     �0�M�H��     ��H�0�L�H��     �T�JH��     �L�����UH��H����H�����I��      L�H��     �T��u
�    �   H��     �T��	vH��     �D    H��     �LH��     ��HT��U�H��     �T�JH��     �L0H��     ��H��D�    �E�����UH����H�����I�/�      L�H��     �D    H��     �    H��     �D    �]���UH��AWSH��0��H�����I�П      L�H�}�H�u�H�E�H�E�H�Eȋ@��-�   �E�H�Eȋ@���2�E��E�,  �E�d   �EԍH��E؍P��E܍p�E���H�}�I��A�  ��I��H�*������H��ЋEԍH��E؍P��E܍p�E���H�}�I��A�������I��H��+������H���H�}ȋMԋU؋u܋E�I��A�������I��H��+������H���H�E�H�HH�E܍P�E���
H���u�I��A�    �������H�S�������H�<I��H�{0������H���H���E��E��m��m�J�EԍH��E؍P��E܍p�E���H�}�I��A�������I��H�*������H��ЋEԍH��E؍P��E܍p�E���H�}�I��A�������I��H��+������H���H�}ȋMԋU؋u܋E�I��A�������I��H��+������H����E�    I�߸    H�x�������H���f�E�f�}�
��   f�}� tl�}� ~ff�}�u_�m�f�E�  H�E�H�xH�E܍P�E��H�E����4�E�H���u�I��A������    ��I��H�6-������H���H��H�m��of�}� �\���H�E�H�xH�E܍P�E��H�E����4�E�H���u�I��A������    ��I��H�6-������H���H���E�H�E�H�PH�U��U҈������H�E��  ��H�Eȋ ��u�H�Eȋ �PH�EȉH�E�H��I��H��\������H���H�E��     �    H�e�[A_]���UH��AWSH��0��H�����I�d�      L�H�}��E���� �E�``` �E���� H�Eȋ@0��(�E�H�Eȋ@,��d�E��E�d   �E�2   �E؍P��E��xH�MȋE�I��A�    �   ��I��H��+������H��ЋE؍P��E܍p�E���H�}ȋM�I��A�ȹ   ��I��H��+������H��ЋE؍P��E܍p�E���H�}ȋM�I��A�ȹ   ��I��H��+������H��ЋEԍP��E܍pH�MȋE�I��A�    �Ѻ   ��I��H��+������H��ЋEԍP��E܍p�E���H�}ȋM�I��A�ȉѺ   ��I��H��+������H��ЋEԍP��E܍p�E���H�}ȋM�I��A�ȉѺ   ��I��H��+������H��ЋEԍP��E܍p�M��E�ȃ�H�}ȋM�I��A�ȉѺ   ��I��H��+������H��ЋEԍP��E܍p�M��E�ȃ�H�}ȋM�I��A�ȉѺ   ��I��H��+������H��ЋEԍP��E܍p�M��E�ȃ�H�M�I��A�    �Ѻ   ��I��H��+������H��ЋE؍P��M܋E�ȍp��E���H�}ȋM�I��A�ȹ   ��I��H��+������H��ЋE؍P��M܋E�ȍp��E���H�}ȋM�I��A�ȹ   ��I��H��+������H��ЋE؍P��M܋E�ȍp��E���H�M�I��A�    �   ��I��H��+������H��АH��0[A_]���UH��AWSH��0��H�����I�.�      Lۉ}܉u؉UԉM�D�E�D�M�H�} u
�    ��  �H   I��H���������H���H�E�H�}� u
�    ��  H�E�H   �    H��I��H�q������H���H�UH�E�H�P@H�E�U�PH�E�P0�E��H�E�PH�E�P,�E��H�E�PH�E��    H�E�P(�E�9�wH�E�P(H�E�P�
�U�H�E�PH�E�P$�E�9�wH�E�P$H�E�P�
�U�H�E�P�U�H�E�P�U�H�E�P H�E��@0    H�E�@0��I��H���������H���H��H�E�H�P8H�E�H�@8H��t.H�E�@0H�U�H�R8H�щ¾    H��I��H�q������H���H�E�@ ��H�E�@��H�E�@��H�E�@��H�E�@L�MA����I��H�*������H���H�E�@��H�E�@��H�E�@��H�E�@L�MA�������I��H��+������H���H�E�H��0[A_]���UH��AWSH��0��H�����I��      L�H�}�H�}� u
������,  I�߸    H�x�������H��҉E�}���   I�߸    H�x�������H��҉E�}�[uqI�߸    H�x�������H��҉E�}�At�}�Bt �2H�Eȋ@,��t&H�Eȋ@,�P�H�EȉP,�H�Eȋ@,�PH�EȉP,��H�E�H��H�xj������H��и    �pH�E�H��I��H�Z�������H���H�E�H�EȋP(H�E�� 9�s=H�E�� ��H�EȉP(H�Eȋ@(��:vH�E��@(    H�E�H��H�xj������H��и    H��0[A_]���UH��AWSH��@��H�����I�y�      L�H�}�H�E�H�@@H�E�H�E�H�@8H�E�H�E�@   H��H�l�������H�<I��H��
������H��ЉE��E�    H�E��@���E���H�EЋ ��u�H�EЋ �PH�EЉ�E�    �!  H�E��@�E�H�E��@ �E�H�E��P,�E�9�u�E�i� �E�����H�E��@��A��H�E��@�U���Ѓ���H�E��@����H�UЋE�I��A���   D��I��H�*������H��ЋE�;E���  H�E�H��H�hm������H���H�E�H�xH�u؋U�H�E��@�M���ȃ�A��H�E��H�E�ȃ�A��H�E�H���u�I��A����D��D��H��I��H�{0������H���H��H�E��@��E�ЉE�H�E�H�xH�u؋E�H�U��R�M���ʃ�A��H�U��J�U�ʃ�A��H���u�I��A����D��D��H�p       H�<I��H�{0������H���H��H�E��@���E�ЉE�H�E�H�xH�u؋E�H�U��R�M���ʃ�A��H�U��J�U�ʃ�A��H���u�I��A����D��D��H��       H�<I��H�{0������H���H���E�    H�m考E��E�;E������H�E��     �H�e�[A_]���UH��AWSH��@��H�����I���      L�H�}�H�E��@b���� ����  H�o�������H�H�t�������H�4H��       H�<I�߸    H�	�������H���H�E��@o��H��x�H*��H��H���H	��H*��X��E�H�����������E��E�    H�E��@o=���?v�E�   H�����������E��)H�E��@o=�� v�E�   H�����������E��E��^E��E�H�E�fHn�H�w�������H�4H�p       H�<I�߸   H�	�������H���H�p       H�<I��H�vv������H��ЉE̋ẺE��H�p       �E�H�H�� �E��}�~�H�        �E�H�H�H��H�w       H�H�t�������H�4H��I�߸    H�	�������H����   H�{�������H�H�t�������H�4H��       H�<I�߸    H�	�������H���H�{�������H�H�t�������H�4H�p       H�<I�߸    H�	�������H��ѐH��@[A_]���UH��H��8��H�����I���      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �CH�E�H�PH�U�� ���E�H�E�H�PH�U�� ���E�E�+E�E�}� u�}� t
�m��}� u��E�����UH��H��8��H�����I�c�      L�H�}�H�uЉŰẺE�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M����E��P��U���u�H�E�����UH��H�� ��H�����I��      L�H�}���U��E�E��E�H�E�H�E��H�E�H�PH�U��U��m��}� u�H�E�����UH��AWSH��0��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E��E�    H�E�H�PH�U�� ����I��H��������H��ЉE�H�E�H�PH�U�� ����I��H��������H��ЉEԋE�+EԉE܃}� u�}� t뗋E�H��0[A_]���UH��AWSH����H�����I�̍      L�H�}�H�u�H�E�H��I��H�vv������H��Љ�H�E�H�H�E�H��H��I��H��s������H���H�E�H��[A_]���UH��H�� ��H�����I�U�      L�H�}�u�H�E�H�E��H�E�� ��9E�uH�E��H�E�H�E�� ��u۸    ����UH��H�� ��H�����I��      L�H�}�H�u�H�E�H�E�H�E�H�E��3H�E��H�E�� 8�u!H�E�� ��H�E�� ��Ѕ�u�    �'H�E�H�PH�U��H�E�H�PH�U�� 8�t����������UH��H��0��H�����I�Z�      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E��  H�E�����UH��AWH��(��H�����I�݋      L�H�}؉uԋU��҉Uԃ}� uOH�U�H��I��H�vv������H��҉�H�E�H���   H�E�� ��tH�E�� ��9E�u	H�E��   H�E�H�E؃�H��űE�i��E�H�E�H�E��H�E�H�E� ������H�E� ��!�%������u%H�E� 3E䍐����H�E� 3E���!�%������t�H�E�H�E��H�E�H�E�� ��tH�E�� ��9E�u�H�E�H��(A_]���UH��H��@��H�����I���      L�H�}�H�u�H�U�H�U�H�U������   H�U�H�������   H�E�    H�E�    H�E�    H�E�    �H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�t�H�E�H+E��'H�U����H�Uȉ�H��H�t������H���H+E�����UH��H����H�����I�~�      L�H�}�H�E�H�E��H�E�H�E�� ��u�H�E�H+E�����UH��AWSH��@��H�����I�/�      L�H�}�H�u��U�H�E�H�E�H�E�H�E��E�    �kH�E�H�PH�U�� ����I��H��������H��ЉE�H�E�H�PH�U�� ����I��H��������H��ЉEԋE�+EԉE܃}� u�}� t
�m��}� u��E�H��@[A_]���UH��H��(��H�����I�j�      L�H�}�H�u��U�H�E�H�E�H�E�H�E��}� u)������2H�E�H�PH�U��H�E�H�PH�U�� 8�u�m��}� u����E�����UH��H��8��H�����I��      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �!H�U�H�BH�E�H�E�H�HH�M����E��E�9E�w�H�E��  �E�����UH��AWH����H�����I�k�      L�H�}�H�u�H�M�H�U�H��H��I��H�@u������H��҉�HE�H�E�� ��tH�E���    H��A_]���UH��AWH��(��H�����I���      L�H�}؉u�H�U�H��I��H�vv������H��҉E��U�H�E�H�H�E��E�    �H�E�� ��9E�uH�E��H�m��E��E�9E�wڸ    H��(A_]���UH��H��0��H�����I�h�      L�H�}�H�u�H�E�H� H�E�H�}� u�    �vH�E�H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u,�}� u
H�E�    �H�E�H���  H�E�H�U�H�H�E���}� u������UH��H��@��H�����I���      L�H�}�H�u�H�E�H�E�H�E�    H�E�    H�E�    H�E�    H�E�� ��u
�    ��   H�E�H��� ��u+�H�E�H�E��H�E�� 8�t�H�E�H+E��   H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�u�H�E�H+E�����UH��H��8��H�����I�x�      L�H�}�H�u�H�U�H�}� uH�E�H� H�E�H�}� u
�    ��   �H�E�H�PH�U�� ���E�H�E�H�E��
�E�;E�u��H�E�H�PH�U�� ���E��}� uۃ}� uH�E�H�     �    �   H�E�H��H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u4�}� u
H�E�    �H�E�H��H�E�H�E��  H�E�H�U�H�H�E���}� u������UH��H����H�����I�A�      L�H�}�H�u�H�u�H�M�H��       H�H��H�|{������H�������UH��AWSH�� ��H�����I��      L�H�}�H�u�H�E�H��I��H�vv������H��ЉE��2�U�H�M�H�E�H��H��I��H��o������H��Ѕ�uH�E��H�E�H�E�� ��uø    H�� [A_]���UH��AWSH�� ��H�����I�O�      L�H�}�H�E�H��I��H�vv������H��Ѓ��E�E��I��H���������H���H�E�H�}� u�    �$�U�H�M�H�E�H��H��I��H��p������H��АH�� [A_]���UH��H��8��H�����I���      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��U�H�E�H�H�E�H�E�H;E�v[H�E�H;E�sQH�E�H�E��E�HE��H�m�H�m�H�E��H�E��H�E�H;E�u��'H�U�H�BH�E�H�E�H�HH�M���H�E�H;E�u�H�E�����UH��AWH����H�����I��      L�H�}�H�u�H�M�H�U�H��H��I��H� s������H���H��A_]���UH��AWH����H�����I���      Lډ}�H���������H�<I�׸    H�ҟ������H�������UH��H����H�����I�J�      L؉}��U���H���������H�Hc��������t�E� �E�����UH��H����H�����I��      L؉}��U���H���������H�Hc��������t�m� �E�����UH��AWSH��0��H�����I��      L�H�}ȉuĉU��M��U�H�E�H��H���������H�<I�߸    I�ҟ������I�A��H�E�H��I��H�Z�������H���H�E�H�E� �E�H�E� 9E�u��H��0[A_]���UH��AWSH�� ��H�����I��~      L�H�}�H�u�H�E�� ��u�    �LH�E�� <wuH�E�H��I��H�d�������H���H�U�H�E�H��H��I��H���������H���H�E�H�E�H�� [A_]���UH��AWH����H�����I�f~      L�H�}�H�U�H��I��H� �������H���H��A_]���UH��AWH����H�����I�~      L�H�}�H�U�H��I��H�9�������H���H��A_]���UH��AWH����H�����I��}      L؉}�H�u�H�M��U�H�Ή�I��H���������H���H��A_]���UH��AWSH�� ��H�����I�|}      L�H�}�H�}� u������VH�E�H��I��H���������H��ЉE�H�E؋@��u+H���������H�H��E�H�։�I��H���������H��ЋE�H�� [A_]���UH��AWH����H�����I��|      L؉}�H�u�H�M��U�H�Ή�I��H�"�������H���H��A_]���UH��AWH����H�����I��|      L�H�}�H�U�H��I��H�u�������H���H��A_]���UH��AWSH��@��H�����I�F|      L�H�}ȉu�H�U�H�}� u	H�E��  H�E�H�E�H�E�H�E��E�    H�E�H��I��H���������H��ЉEԃ}����   H�E��@��u7�}�u�}� ~+H���������H�H��E�H�։�I��H���������H��Ѓ}�
tk�E�;E�}E�}�u�}� ~H�E�H;E�vH�m��m��:�}��^���H�E�H�PH�U�UԈ�E��D����}�u�}� ~�m���E��)�������}�~	H�E��  ��Eԉ�H�E�H�E�H��@[A_]���UH��AWSH�� ��H�����I��z      L�H�}�H�u�H�}� u�    �^�E�    �2�E�Hc�H�E�H�� ��H�U�H�։�I��H�"�������H��ЃE�H�E�H��I��H�vv������H��ЋU�9�w��E�H�� [A_]���UH��AWH��(��H�����I�Hz      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I�}�������I�A��H��(A_]���UH��AWH��(��H�����I��y      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I�>�������I�A��H��(A_]���UH��AWH����H�����I��y      L�H�}�H�U�H��I��H�f������H���H��A_]���UH��AWH����H�����I�Cy      L�H�}�H�U�H��I��H��������H��ҐH��A_]���UH��AWH��(��H�����I��x      L�H�}�H�u��U܋U�H�u�H�M�H��I��H���������H���H��(A_]���UH��H����H�����I��x      L�H�}�H�}� u������!H�E��P#H�E���+  9�r�������    ����UH��AWH����H�����I�Ex      L�H�}�H�U�H��I��H���������H���H��A_]���UH��AWSH��`  ��H�����I��w      L�H������H������H�������E�    �E�    �  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H���������H���	E�}���  �E�H��    H��k  H�H��k  H�>��H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E��E�H������H�։�I��H��������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�}� t(H������H�E�H��H��I��H��������H����O  H������H��H���������H�<I��H��������H����   H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E�H�������E�H�։�I��H�˯������H���H������H������H��H��I��H��������H����w  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������
   H��H��I��H�E�������H���H������H������H��H��I��H��������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������   H��H��I��H��������H���H������H������H��H��I��H��������H����  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�EȾ   H��fHn�I��H� �������H���H������H������H��H��I��H��������H����]  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eк
   H��H��I��H���������H���H������H������H��H��I��H��������H����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ
   H��H��I��H�E�������H���H������H������H��H��I��H��������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ   H��H��I��H�E�������H���H������H������H��H��I��H��������H����G  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�E�   H��fHn�I��H� �������H���H������H������H��H��I��H��������H����   H������H�ƿ%   I��H��������H��ЋE�Hc�H������H�� ��H������H�։�I��H��������H����4�E�Hc�H������H�� ��H������H�։�I��H��������H��ЃE��E�Hc�H������H�� ��������    H��`  [A_]���UH��H����H�����I�ko      L؉��E��E�    �E��S��%wa��H��    H��d  H�H��d  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��n      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��H�� ��H�����I��m      L�H�}�H�u�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E�����UH��AWSH��  ��H�����I�dm      L�H������H������H��x����E�    H������H�E�f�E�  �E� �E�    �/  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H�_�������H���	E܃}���  �E�H��    H�Bc  H�H�7c  H�>��H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E��E�H�U�H�E�H��H��H��������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H�}� t'H�U�H�E�H��H��H��������H���H�E��e  H�E�H���������H�4H��H��������H���H�E��7  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E�H�������E�H�։�I��H�˯������H���H������H�E�H��H��H��������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������
   H��H��I��H�E�������H���H������H�E�H��H��H��������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������   H��H��I��H��������H���H������H�E�H��H��H��������H���H�E��3  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�E��   H��fHn�I��H� �������H���H������H�E�H��H��H��������H���H�E��x  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�E��
   H��H��I��H���������H���H������H�E�H��H��H��������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ
   H��H��I��H�E�������H���H������H�E�H��H��H��������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ   H��H��I��H�E�������H���H������H�E�H��H��H��������H���H�E��e  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�Eо   H��fHn�I��H� �������H���H������H�E�H��H��H��������H���H�E��   H�E�H���������H�4H��H��������H���H�E�fǅ����  �E�Hc�H������H�� ������H������H�E�H��H��H��������H���H�E��8�E�Hc�H������H�� �E�H�U�H�E�H��H��H��������H���H�E��E��E�Hc�H������H�� �������H�E��  H�U�H������H)�H��H�Ā  [A_]���UH��H����H�����I��d      L؉��E��E�    �E��S��%wa��H��    H��[  H�H��[  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��c      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H���������L��Љ�<�����<���Hc�H�����H��  ��<���H���   A_]���UH��AWH���   ��L�����I��b      M�H����������H�����H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H����������H�����H��M��H���������L��Љ�<�����<���H���   A_]���UH��AWSH��0��H�����I��a      L�H�}؉u�H�U�H�M��}�   v
�    �   H�U�H�E�H��H��       H�<I��H���������H��ЉE�}���  ~�   �I�E�E�}� ~:�U�H�E�H��       H�4H��I��H��p������H��ЋE�Hc�H�E�H��  �E�H��0[A_]���UH��AWH����H�����I�"a      L؉}�H���������H�H�
�U�H�Ή�I��H�"�������H���H��A_]���UH��AWSH�� ��H�����I��`      L�H�}�H�}� tj�E�    �?H���������H�H��E�Hc�H�E�H�� ��H�։�I��H�"�������H��ЃE�H�E�H��I��H�vv������H��ЋU�9�w���H�� [A_]���UH��AWH���   ��L�����I�`      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I�(_      M�H��8���H��0���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�H���������I�<M�׸    H�ҟ������L�������UH��AWH����H�����I��^      L�H�}�H�U�H��I��H�,�������H��ҐH��A_]���UH��AWH��(��H�����I�>^      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H���������H��Ѹ    H��(A_]���UH��AWH��(��H�����I��]      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H���������H����H�E�H�E�� < tH�E�H   H9E�sH�E�� <
u�H�E��  H�E�H;E�����H��(A_]���UH��AWSH��0��H�����I�6]      L�H�}�H�uЉỦM�H��      H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H���������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H��      H�H�E�H��      �0H��      �D �}�u-�U�H�E�    H��I��H�z�������H���H�U�H��   �}�u+�U�H�E�    H��I��H���������H��Љ�H�EЉ�[�}�u,�U�H�E�    H��I��H���������H��Љ�H�E�f��)�U�H�E�    H��I��H���������H��Љ�H�EЈ�    H��0[A_]���UH��AWSH��0��H�����I��[      L�H�}�H�uЉỦM�H��     H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H���������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H��     H�H�E�H��     �0H��     �D �}�u'H�E�H��I��H���������H����Z�H�E�� �+�}�u%H�E�H��I��H���������H���fH~�H�U�H��    H��0[A_]���UH��SH��8��H�����I�WZ      L�H�}�H�u�H�U��E�    �E�    ��  �E�    �E�Hc�H�E�H�� ������%��  �E��E�Hc�H�E�H�� ������lu�E��E�   �E�Hc�H�E�H�� ����H���������H���	E�}��o  �E�H��    H�dR  H�H�YR  H�>��H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H���������H�����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H��������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�_�������H����?  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H�����   H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H����jH�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�_�������H������E��E�Hc�H�E�H�� ��������E�H��8[]���UH��H����H�����I��U      L؉��E��E�    �E��S��%wa��H��    H�SO  H�H�HO  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I�MU      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I�bT      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��H����H�����I�rS      L؉}�H�u�H�}� u������w�}��u������jH�E��@#��tH�E��@#�P�H�E��P#H�E��@#H�U��J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U���E�����UH��AWSH����H�����I��R      L�H���������H�H� H��I��H���������H��ЉE�}��t+H���������H�H��E�H�։�I��H���������H��ЋE�H��[A_]���UH��AWH��(��H�����I�1R      L�H�}�H�u�H�U�H���������H�<I�ϸ    H�ҟ������H�������UH��H����H�����I��Q      L�H�}��	   H�E�H���r�����UH��SH����H�����I��Q      L�H�}�H�}� u.H��     H�<H��������H���H��     H��H�E�H��H��������H���H�E�H��[]���UH��AWSH��0��H�����I�Q      L�H�}�H�u�H�E�H���������H�4H��I��H���������H���H�E�H�}� u
������   �E�    H�E�H��I��H�vv������H��ЉE܃}�`~	�E�   �$H�E�H�P+H�E�H��H��I��H��s������H���H�E��@���H�E��PH�E�H��I��H���������H��ЋE�H��0[A_]���UH��H��0��H�����I�)P      L؉}�H�u�H�E�H�E��E܉E��E�    �}� y,H�E�H�PH�U�� -�}�   �u�E�����E���E��؉E�H�E�H�E�M�Hc�Hi�gfffH�� ��������)�����)��ʉЍH0H�E�H�PH�U�ʈ�E�Hc�Hi�gfffH�� ����)ЉE�}� u��}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWSH��@��H�����I��N      L�H�}�H�u��U�H�}� u#H�E�H�E�H�E�H�PH�U�� 0H�E��  �  H�E�H�E؋E�Hc�H�E�H�H�E��3H�E؃��E�H�m��}�	~�7   ��0   �U��H�m���H�E�H�E�H;E�wËE�Hc�H�E�H��  H�E�H�E��E�    �8H�E�� <0uH�E��"H�U�H�E�H��H��I��H��s������H�����E��E�;E�|�H�E�H�E�H�E�H��I��H�vv������H��Љ�H�E؋E�H�U�)Љ�H�M�H�E�HȾ    H��I��H�q������H���H��@[A_]���UH��AWH����H�����I�kM      L؉}�U�    ��I��H��������H���H��A_]���UH��AWH����H�����I�M      L؉}�u�U��U��I��H���������H���H��A_]���UH��AWH����H�����I��L      L�H�}�H�U�H��I��H�������H��ҐH��A_]���UH��AWH����H�����I��L      L�H�}�u�M�H�U��H��I��H�������H���H��A_]���UH��H����H�����I�2L      L؉}�u�E��}�E��E��}�ЉE��}� x�E���y�E����E��E�+E�E��!�}� y�E���~�E����E��U��E�ЉE�H�E�����UH��H�� ��H�����I��K      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H�� ��H�����I� K      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H��H��H�����I�VJ      L�H�}�H�u��U�H�E�H�E�H�E�H�PH�U�� ���E�E���H���������H�H������ ��uǃ}�-u�E�   H�E�H�PH�U�� ���E��"�E�    �}�+uH�E�H�PH�U�� ���E�}� t�}�u9�}�0u3H�E�� <xtH�E�� <XuH�E�H��� ���E�H�E��E�   �}� u�}�0u�   ��
   �E��}� t	H��   ������H�E�E�Hc�H�E�H�H��H�ЉE؋E�Hc�H�E�H�H��H�E�}� t�}� ~�E�)E�H�E��]�H�E�    �E�    �E���H���������H�H��������t�m�0�[�E���H���������H�H���������5  �E���H���������H�H��������t�7   ��W   )E�E�;E���   �}� ��   �}� tgH�E�H;E�|H�E�H;E�u0�E�;E�~(�E�����H�E�   �H���������H�� �����   �E�   �E�H�H�U�H��H�E��E�H�H)E��eH�E�H;E�H�E�H;E�u-�E�;E�~%�E�����H�E����H���������H�� �����$�E�   �E�H�H�U�H��H�E��E�H�HE���H�E�H�PH�U�� ���E��y������H�}� t�}� t
H�E�H���H�E�H�U�H�H�E�����UH��AWH����H�����I�"G      L�H�}�H�M�
   �    H��I��H���������H���H��A_]���UH��AWH����H�����I��F      L�H�}�H�M�
   �    H��I��H���������H���H��A_]���UH��AWAVAUATSH����H�����I�qF      L�H�}�H�uȉU�L�eп    L��L�`� �؉���H���������H�H������ ��uЃ�-u�   L��L�`� �����+uL��L�`� �؃}� t�}�u-��0u(A�$<xt	A�$<XuI�D$� ��I���E�   �}� u��0u�   ��
   �EċE�Hc������    H��I�ǋE�Hc������    H��H�Љ�A�    A�    ����H���������H�H��������t��0�T����H���������H�H��������tz����H���������H�H��������t�7   ��W   )�;]�}GE��x
M9�wM9�u��9�~A������A�   �E�H�L��Hc�I�L��L�`� ���;������E��yA�����H���������H�� "   �	����tI��H�}� tE��tI�D$��H�E�H�U�H�L��H��[A\A]A^A_]���UH��H����H�����I�.D      L؉}��   �   ���r����UH��AWSH����H�����I��C      L�H�}�H�E�H���������H�4H��I��H� s������H��Ѕ�uH���������H�H� ��    H��[A_]���UH��AUATSH�� ��H�����I�{C      L�H�}�H�u�H�8     ��E�L�e�H�]�E�,$L��L�`��H��H�XD�(�m��}� uې�H�� [A\A]]���UH��H��8��H�����I�C      L�H�}�H�u�H�U�H�8     ��E�H�E�H�E�H�E�H�E�H�E�H�E�H�E�� ���E�H�E�H�PH�U�H�U���H�E�H�PH�U�H�U���H�E�H�PH�U��U���m��}� u�������UH��SH��H��H�����I�VB      L�H�}�H�u�H�8     ��E�H�E�H+E��EȋE�9E���  �E�����EȺ    ��E��EȋU�H�E�H�H�E�H�E�H�E�H�E�H�E�E�H�H��H��H�E�H�H�E�H�E�H;E�sjH�0     H�H�U�H�E�H��H���щEă}� u/�E�H�H��HE�H�U�H�E�H��H��H�t�������H�����  �}� y�E�H�HE���  �H�E�H;E���   H�0     H�H�U�H�E�H��H���щEă}� u)�E�H�HE�H�U�H�E�H��H��H�t�������H���뢃}� ��   H�E�H;E�uA�E�H�HE�H�U�H�M�H�E�H��H��H��������H��ЋE�H�HE�H�E�H�E��M���H�U�H�E�H��H��H�t�������H��ЋE�H�H��HE��E�H�HE���   �E�H�H��HE�����H�E�H;E���   H�E�H+E�H��H�E�H+E�H9�|4�E�Hc�H�E�H�H�E�H��H��H���������H���H�E�H�E������H�U�H�E�H��H��H���������H��ЋE�Hc�H�E�H�H�E������E�H�H��HE�H�U�H�M�H�E�H��H��H��������H��ЋE�H�H��HE�H�E�H�E������H��H[]���UH��H�� ��H�����I�e?      L�H�}��u�U�H�M�H�0     H�U�H��U�H�8     ��U��U���H�U�H�H�U�H��H��H���������H��А����UH��AWH����H�����I��>      L�H�}�H���������H�<I�׸    H�ҟ������H��Ѹ����H��A_]���UH��H��@��H�����I��>      L�H�}�H�u�H�U�H�U��H�E�H�U����H���������H�Hc���҃� ��u��E�    H�U���҃�+t��-u�E�   H�E�H� ���������E��E�    �E�    �E�    �;�M�H����������Y�H�U���҃�0�*��X��E�H�E��E�H�U����H���������H�Hc���҃���u�H�U����.uuH�E��?�M�H����������Y�H�U���҃�0�*��X��E�H�E��E��E�H�U����H���������H�Hc���҃���u��U�)U�}� uH� �������f���  �}� t�E�H��������f(fW��E�H�U����etH�U����E��   �E�    H�E�H�U���҃�+t��-u�E�   H�E��E�    �%�M܉����҉�H�U���҃�0ʉU�H�E�H�U����H���������H�Hc���҃���u��}� t�U�)U���U�U�}����|	�}�   ~H�����������   H����������E��E�E܃}� yF�]��A�E܃���t&�}� y�E��^E��E���E��YE��E��}��E��Y��E��}� u�H�}� tH�E�H�U�H��E�����UH��H����H�����I�S;      L؉}�H�E�   �E�    �H�U�H��H��H�H�H�E��E��E�;E�|�H�E�����UH��AWSH��@��H�����I��:      L��E�H�}��u�H�}� u	H�E��  H�E�H�E�H�(�������f��f/E�v,H�E�H�PH�U�� -�E�H�0�������f(fW��E��E�H�@�������f/s�E��H,�H�E��/�E�H�@���������\��H,�H�E�H�       �H1E�H�E�H�E�H�E�H��x�H*��H��H���H	��H*��X��M��\�f(��EȋE���H���������H���H��x�H*��H��H���H	��H*��X��YE�H�@�������f/s�H,�H�E��*H�@���������\��H,�H�E�H�       �H1E�H�E�H�E�H�M�H�U�H�E�H� �������H�43H��I�߸    I�	�������I�A��H�E�H��@[A_]���UH��AWH����H�����I�9      L�H�}�H�U�    H��I��H�l�������H���H��A_]���UH��AWH����H�����I��8      L�H�}�H�u�H�M�H�U�H��H��I��H�l�������H����Z�H��A_]���UH��AWH��(��H�����I�]8      L�H�}�H�u�H�M�H�U�H��H��I��H�l�������H����E��E�H��(A_]���UH��H����H�����I�8      L؉}��E����3E�)�����UH��H��@��H�����I��7      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�    H�}� y>H�E�H�PH�U�� -H�       �H9E�uH��������H�E�H�E��H�E�H��H�E�H�E�H�E�H�M�H�gfffffffH��H��H��H��H��?H)�H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U��ʈH�M�H�gfffffffH��H��H��H��H��?H)�H��H�E�H�}� u�H�}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U߈H�E�H;E�w�H�E�����UH��AWH��8��H�����I�U6      L�H�}�H�uЉU�H�U�H�U�H�}� yH�U�H�JH�M��-H�]�H�U�H�U��}�u$H�M�H�u�   H��I��H��������H����H�M�H�U�H��H��H�'�������H���H�E�H��8A_]���UH��H��0��H�����I��5      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E�H�M�H���������H��H��H��H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U�ʈH�E�H���������H��H��H��H�E�H�}� u�H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWH��8��H�����I��4      L�H�}�H�uЉU�H�U�H�U�H�U�H�U��}�u$H�u�H�M�   H��I��H��������H����H�M�H�U�H��H��H�L�������H���H�E�H��8A_]���UH��H����H�����I�4      L؉}������UH����H�����I��3      Lظ   ]���UH��H����H�����I��3      L�H�}��    ����UH��H����H�����I��3      L�H�}�H���������H�H� ����UH��H����H�����I�_3      L�H�}�H���������H�H� ����UH��H�� ��H�����I�$3      L�H�}��u�H�U�H�M�    ����UH����H�����I��2      Lظ    ]���UH��H����H�����I��2      L��E�H�H�������f������UH��H����H�����I��2      L��E�H�H�������f������UH��H����H�����I�Q2      L��E��}�H�H�������f������UH��H����H�����I�2      L��E�H�}�H�H�������f������UH��H����H�����I��1      L��E��M�H�H�������f������UH��H��(��H�����I��1      L��E��M��E��U��U��E��E��E������������������������������]��E�����UH��H����H�����I�,1      L��E����E����]��E�����UH��H����H�����I��0      L��E�H�P�������f������UH��H����H�����I��0      L��E�H�X�������f������UH��H����H�����I�0      L��E�H�`�������f������UH��H����H�����I�F0      L��E�H�h���������E��E�����UH��H����H�����I�0      L��E�H�p�������f������UH��H����H�����I��/      L��E�H�x�������f������UH��H����H�����I��/      L��E�H���������f������UH��H����H�����I�W/      L��E�H���������f������UH��AWH����H�����I�/      L��E��E�H���������H�f(�fHn�I��H�Z�������H���H��A_]���UH��H����H�����I��.      L؉}�H�u�    ����UH��AWH����H�����I��.      Lډ}�H�u�H���������H�<I�׸    H�ҟ������H�������UH��AWH��(��H�����I�5.      Lى}�H�u�H�U�H���������H�<I�ϸ    H�ҟ������H�������UH��AWSH�� ��H�����I��-      L�H�}�H���������H�<I�߸    H�ҟ������H����E�    �.�E�H�H��    H�E�HЋ ��I��H�О������H��ЃE��}�?~̸����H�� [A_]���UH��AWH����H�����I�B-      L�H�}�u�H���������H�<I�׸    H�ҟ������H�����f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f�                                                                    ~ � � � � � � � � ~             ~ � � � � � � � � ~                 l � � � � | 8                   8 | � | 8                   < < � � �   <                < ~ � � ~   <                      < <              � � � � � � � � � � � � � � � �           < f B B f <           � � � � � � � � � � � � � � � �        2 x � � � � x             < f f f f <  ~               ? 3 ? 0 0 0 0 p � �              c  c c c c g � � �               � < � < �             � � � � � � � � � � �               > � >                  < ~    ~ <                f f f f f f f   f f              � � � {                | � ` 8 l � � l 8  � |                       � � � �              < ~    ~ <  ~              < ~                           ~ <                      �                         0 ` � ` 0                         � � � �                       ( l � l (                      8 8 | | � �                   � � | | 8 8                                                 < < <                  f f f $                             l l � l l l � l l           | � � � |   � � |               � �   0 ` � �             8 l l 8 v � � � � v           0 0 0 `                             0 0 0 0 0 0               0         0                   f < � < f                         ~                                    0                     �                                                           0 ` � �             8 l � � � � � � l 8              8 x       ~             | �    0 ` � � �             | �   <    � |               < l � �                 � � � � �    � |             8 ` � � � � � � � |             � �     0 0 0 0             | � � � | � � � � |             | � � � ~     x                                                       0                  0 ` 0                      ~     ~                     ` 0      0 `             | � �                       | � � � � � � � |              8 l � � � � � � �             � f f f | f f f f �             < f � � � � � � f <             � l f f f f f f l �             � f b h x h ` b f �             � f b h x h ` ` ` �             < f � � � � � � f :             � � � � � � � � � �             <         <                   � � � x             � f f l x x l f f �             � ` ` ` ` ` ` b f �             � � � � � � � � � �             � � � � � � � � � �             | � � � � � � � � |             � f f f | ` ` ` ` �             | � � � � � � � � |           � f f f | l f f f �             | � � ` 8   � � |             ~ ~ Z       <             � � � � � � � � � |             � � � � � � � l 8              � � � � � � � � � l             � � l | 8 8 | l � �             f f f f <     <             � � �   0 ` � � �             < 0 0 0 0 0 0 0 0 <               � � � p 8                 <         <          8 l �                                                   �       0                                     x  | � � � v             � ` ` x l f f f f |                   | � � � � � |                < l � � � � v                   | � � � � � |              6 2 0 x 0 0 0 0 x                   v � � � � � |  � x       � ` ` l v f f f f �                 8      <                        f f <       � ` ` f l x x l f �             8         <                   � � � � � � �                   � f f f f f f                   | � � � � � |                   � f f f f f | ` ` �             v � � � � � |                � v f ` ` ` �                   | � ` 8  � |              0 0 � 0 0 0 0 6                    � � � � � � v                   � � � � � l 8                   � � � � � � l                   � l 8 8 8 l �                   � � � � � � ~   �             � �  0 ` � �                 p                                        p         p                       v �                        8 l � � � �                               ��� ��� ~~~                                 uuu ��� ��� ���                                 ��� ��� ��� ��� ;;;                          ��� ��� ~~~ ��� ���                         ��� ��� ���     ��� ���                         ��� ���      ��� ��� ppp                 @@@ ��� ���         III ��� ���                 ��� ��� ��� ��� ��� ��� ��� ���                 ��� ���                 zzz ��� ���         ``` ��� ���                     ��� ���         ��� ��� MMM                     ��� ��� bbb     ��� ���                         ||| ��� ���      ��CFiles SIM
      Entrada maior que o limite
 Erro ao criar o arquivo "%s"
       Error ao criar o arquivo "%s", atingio o limite de arquivos na entrada de directorio
   Panic: __malloc, sem espaco na tabela de alocacao
      panic: realoc sem espaco, %lx size = %d %d
 PWD BitMAP error
 Not suport BitMAP 4-bit Not suport BitMAP > 8-bit ____ none
 File name    KIB MiB GiB ./ File %s %lf            �@      �A      0Astrerrorr
              (((((�AAAAAABBBBBB                                �Dubug: %s %x %x
        (null)  ��������(���������������i����������������������p�������p�����������������������������������������������������������������������������������������������,�������ޘ��������������B�������B�������`���������������������������������������{���������������������������������������������������������������������������������������W�������i���������������������������������������i�������������������������������������������������������������������������������`���������������r�����������������������{�������(null) %        ��������Ϝ������Z����������������������k�������������������������������������������������������������������������������������������������������������Ԡ��������������6���������������������6�������l�������l�������l�������l�������Q�������l�������l�������l�������l�������l�������l�������l�������l�������l�������l�������-�������?�������l�������c�������Z�������l�������?�������l�������l�������l�������l�������l�������l�������l�������l�������l�������6�������l�������H�������l�������l�������Q�������panic: sscanf()
        �����������������������w����������������������O�������O�������������������������������������������������������������������������������������������������������'�������������������������������ǰ�������������������������������������������������������������������������������������������������������������������������������������а�������������������������������������а������������������������������������������������������������������������������ǰ��������������ٰ�����������������������������panic: freopen()
 r+ PWD call system funtion error. 
                 $@       �        %lu.%lu                �              �C                                                                        �_�
�@panic: signal()
 panic: sigaction()
 panic: setjmp()  panic: longjmp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �C �     �     �   @L �   �C �   �T �   �C �      �   �C �      �   �C �    4 �   �C �   D �                                   �3 �   �3 �   �3 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  zR x�  ,      @����   E�CG����B�A�          L   �����   E�CG��  $   l   v����    E�CG��w�B�A�(   �   ����Z   E�CG��G�B�A�      �   ���   E�C�   �   ����    E�C��       �����    E�C��        ���p    E�CF�`�A�$   D  a����    E�CG����B�A�$   l   ���r    E�CG��_�B�A�(   �  j���   E�CG��	�B�A�   $   �  Z����   E�CF���A�       �  ����    E�CE���A�      �����    E�CE���A�   0  .����    E�C��    P  ����A    E�Cx�      p  ���i    E�C`�        �  R���U    E�CL�    �  ����U    E�CL�    �  ����i    E�C`�    �  ���g    E�C^�      L����    E�C�� $   4  ����   E�CE�{�A�      \  u���9    E�Cp�  $   |  �����    E�CG����B�A�   �  O���^    E�CU� (   �  ����   E�CG���B�A�   (   �  v����   E�CG����B�A�   (     ���]   E�CG��J�B�A�   (   H  E���   E�CG��l�B�A�   (   t  ����D   E�CJ��.�B�A�   (   �  ����:   E�CG��'�B�A�   $   �  ����    E�CG����B�A�   �  �����    E�C��      J����    E�C�� (   4  �����   E�CJ����B�A�   (   `  ����i   E�CG��V�B�A�   (   �  ����H   E�CG��5�B�A�   (   �  ���e   E�CJ��O�B�A�      �  S���a    E�CX�      ����9    E�Cp�      $  �����    E�CF�w�A�(   H  ���'   E�CG���B�A�   $   t  ���   E�CE���A�   $   �  �����   E�CF���A�      �  ^���    E�C��    �  >����    E�C�� (     ���O   E�CG��<�B�A�   $   0  %����    E�CG����B�A�(   X  ����C   E�CG��0�B�A�      �    ��k    E�Cb� $   �  K ���    E�CG����B�A�   �  ���    E�C�� $   �  ���   E�CE��A�   $     n���    E�CG����B�A�$   <  ����    E�CG����B�A�(   d  ����   E�CG����B�A�   (   �  ��j   E�CG��W�B�A�       �  P���    E�CE���� (   �  ���   E�CG���B�A�       	  ����    E�CE���� (   0	  s���   E�CG��q�B�A�   $   \	  ���   E�CG����B�A�   �	  ���9    E�Cp�     �	  ���+    E�Cb�     �	  ����    E�C��     �	  ;���   E�CE����   
  ���I    E�C@�     (
  ��u    E�CE�f�A�(   L
  W���   E�CG����B�A�   (   x
  ���   E�CG����B�A�   $   �
  ����    E�CG����B�A�,   �
  x��2   E�CG���B�A�       (   �
  z��D   E�CG��1�B�A�   $   (  ����    E�CG����B�A�(   P  	���   E�CG����B�A�   ,   |  ���   E�CG����B�A�       ,   �  o!��   E�CG���B�A�       (   �  ]#���   E�CG��s�B�A�   $     �$���    E�CG����B�A�(   0  v%��   E�CG��
�B�A�   $   \  g)���    E�CG����B�A�$   �  �)��   E�CF��A�   (   �  �*���   E�CG����B�A�   $   �  U/���    E�CG����B�A�(      0��5   E�CG��"�B�A�   $   ,  1��k    E�CG��X�B�A�   T  Y1���    E�C��    t  �1���    E�C��    �  �2��X    E�CO� ,   �  �2��l   E�CG��Y�B�A�       ,   �  6��6   E�CG��#�B�A�       (     9��D   E�CG��1�B�A�   (   @  3;��q   E�CG��^�B�A�   (   l  x<���   E�CG����B�A�   (   �  <?���   E�CG����B�A�      �  �A���    E�C��    �  B��w    E�Cn�      pB��b    E�CY� $   $  �B���    E�CG����B�A�$   L  EC��z    E�CG��g�B�A�   t  �C��a    E�CX�    �  �C���    E�C��    �  RD��{    E�Cr� $   �  �D��+   E�CF��A�      �  �E��6   E�C-�     �F��L    E�CC� $   <  �F���    E�CG����B�A�   d  �G���    E�Cw�    �  �G��}    E�Ct� $   �  OH��r    E�CF�b�A�    $   �  �H���    E�CF���A�       �  I���    E�C��      �I��3   E�C*�   4  �J��7   E�C.�   T  �K��W    E�CN� $   t  L���    E�CG����B�A�$   �  rL���    E�CG����B�A�   �  �L���    E�C�� $   �  �M��V    E�CF�F�A�         �M��P    E�CF�       ,  �M��U    E�CL�    L  N��U    E�CL� $   l  TN���    E�CG����B�A�$   �  �N���    E�CG����B�A�$   �  <O��K    E�CF�{�A�     $   �  _O��K    E�CF�{�A�     $     �O��S    E�CF�C�A�    $   4  �O���    E�CG����B�A�$   \  P��S    E�CF�C�A�    $   �  HP��K    E�CF�{�A�     ,   �  kP��[   E�CG��H�B�A�       $   �  �Q���    E�CG����B�A�$     R��]    E�CF�M�A�    $   ,  GR��]    E�CF�M�A�    $   T  |R��K    E�CF�{�A�     $   |  �R��L    E�CF�|�A�     $   �  �R��Y    E�CF�I�A�       �  �R��Y    E�CP� $   �  -S��K    E�CF�{�A�     (     PS���   E�CJ��{�B�A�       @  �[���    E�C��     $   d  ;\���    E�CI���A�       �  �\��l    E�Cc� (   �  J]���   E�CJ����B�A�       �  �e���    E�C��     $   �  yf��   E�CI���A�    $   $  Rg���    E�CI���A�    $   L  h���    E�CG����B�A�$   t  �h��\    E�CF�L�A�    $   �  �h���    E�CG����B�A�$   �  zi���    E�CI���A�       �  Gj���    E�CI�    $     �j��L    E�CF�|�A�         4  �j��e    E�CF�U�A�    X  -k���    E�CF���A�(   |  �k���   E�CG����B�A�   (   �  #m��=   E�CG��*�B�A�   $   �  4n��\   E�CE�M�A�      �  hr���    E�C�� $     �r���    E�CI���A�    $   D  �s���    E�CI���A�       l  �t���    E�C�� $   �  u���    E�CG��z�B�A�   �  yu��Y    E�CF�       �  �u��9    E�Cp�  $   �  �u���    E�CE�q�A�    $     #v���    E�CG����B�A�   D  �v��G   E�C>�,   d  x��u   E�CG��b�B�A�       $   �  _y��M    E�CF�}�A�     $   �  �y��O    E�CF��A�     $   �  �y��L    E�CF�|�A�     $     �y��S    E�CF�C�A�       4  �y���    E�C�    T  bz���    E�C��    t  �z���    E�C��    �  v{��2   E�C)�$   �  �~��U    E�CF�E�A�    $   �  �~��U    E�CF�E�A�    4     �~��L   E�CM�����-�B�B�B�B�A�      <  ����7    E�C       $   \  ���w    E�CG��d�B�A�(   �  \���{    E�CI���d�B�B�A�   �  �����    E�C�� $   �  9����   E�CE���A�       �  ����    E�Cx�     $     `���\    E�CF�L�A�       D  ����5   E�C,�   d  ����_    E�CV� ,   �  ����   E�CG����B�A�       $   �  ����P    E�CF�@�A�    $   �  ˊ��Z    E�CF�J�A�    $     ����^    E�CF�N�A�       ,  3���4    E�Ck�     L  G���v   E�Cm�$   l  �����    E�CF���A�       �  $����    E�C�� $   �  �����    E�CF���A�       �  j���*    E�Ca�     �  t���'    E�C^�       {���/    E�Cf�     <  ����;    E�Cr�     \  ����;    E�Cr�     |  ����:    E�Cq�     �  ڎ��'    E�C^�     �  ���9    E�Cp�     �  ����9    E�Cp�     �  ���<    E�Cs�       /���=    E�Ct�     <  L���>    E�Cu�     \  j���n    E�Ce�    |  ����;    E�Cr�     �  ӏ��9    E�Cp�     �  ���9    E�Cp�     �  ���9    E�Cp�     �  ���D    E�C{�        B���9    E�Cp�     <   [���9    E�Cp�     \   t���9    E�Cp�     |   ����9    E�Cp�  $   �   ����a    E�CF�Q�A�       �   ߐ��2    E�Ci�     �   ���T    E�CF�    !  )���X    E�CF�$   !  e����    E�CG����B�A�   D!  ؑ��T    E�CF�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    GCC: (Ubuntu 9.3.0-17ubuntu1~20.04) 9.3.0                                        �                    �                  @ �                 p@ �                 �@ �                 �@ �                  ` �                                     ��                     ��_ cole _             ��                )        �           X         �           0    ��                7    ��                A      h2 �           F      n2 �           K    ��                R    ��                A      x2 �           F      �2 �           X      �2 �           �   ��                ]     �@ �          A      3 �           F      H3 �           m    ��                t    ��                A      t3 �           {    ��                �    ��                �    ��                �    ��                A      x3 �           F      �3 �           X      �3 �           �    ��                �    ��                �    ��                �     �  �         �    ��                �    ��                A      �3 �           �    ��                �     �@ �          �    �@ �          �     �@ �          A      �3 �           �    ��                �    ��                A      �3 �           �    ��                   ��                    �@ �                A �                �@ �          �     �  �   �      -    ح  �   �      2     �3 �           7     �3 �           <     �3 �           A     �3 �           F     �3 �           K      4 �           P     �3 �           U     �3 �           [   ��                d   ��                m   ��                v   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                   ��                   ��                     A �             ��                '   ��                0   ��                :   ��                D   ��                A      4 �           O   ��                W   ��                a   ��                k   ��                A       5 �           s   ��                {   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �    ��  �   �       A      85 �           �   ��                �   ��                �    ��  �   �       A      07 �           F      77 �           �   ��                   ��                    ��                    @A �             ��                �   ��                �   ��                   ��                A      09 �           &   ��                /   ��                9    $�  �   e       p    ��  �   �       N    +�  �   �      C    @A �          M    ��  �   =      T    @B �          �    h�  �   �       0   ��                1   ��                ^   ��                g   ��                q   ��                A      8; �           {   ��                �    @C �   `       �   ��                A      J; �           �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                A      M; �               ��                    �C �              �C �              ��  �   {           _�  �   �            �  �   �      $   ��                A      Q; �           -   ��                A      p; �           F      x; �           X      �; �           6   ��                =     �   _       A      �; �           F      �; �           X      �; �           2     �; �           H   ��                O   ��                X   ��                b   ��                h   ��                o   ��                v   ��                w   ��                ~   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                A      �; �           �   ��                �   ��                �   ��                A      �; �           �   ��                A      �; �           �   ��                A      �; �           �   ��                A      �; �           �   ��                A      �; �           �   ��                A      �; �           �   ��                A      �; �           �   ��                A      �; �           �   ��                A       < �           �   ��                �   ��                A      < �           F      < �           �   ��                A      -< �           F      >< �                ��                    p@ �                 �   T       %    U6  �         �    @�  �   \       8    ��  �         B    o  �   �       M    
�  �   {       T    � �   9       X    8 �   ;       ]    � �   �       d    l�  �   �       h    5  �   �       x    �  �   7      T    B�  �   �       �    �C �          �    ��  �   �      �    ��  �   �       �      �               �j  �   �       �      �           �    ʿ  �   P       �    �
 �   �           D �          �    @L �          �    ��  �   �       �    z�  �   �       �    �C �          �    �_  �   �      �    ��  �   U       �    2{  �   u       �    m�  �   w       �     �   9       �    �T �          �    � �   9       �     �   ^           `2 �              �#  �   �           �  �   �       E    �  �   �           �  �   [      "    TG  �   :      .    �I  �   �       >    w�  �   q      ~
    ��  �   �       J    �  �   w            =�  �   �      Q    �w  �   �       `    �~  �   �      h    ��  �   L       o    � �   v      �    ��  �   �       v    �  �   U       ~    � �   \       �    ��  �   Y       �    ��  �   M       �    ��  �   K        
    �C �          �     D �          �    u�  �   �       �    #x  �   �      �     �   <       �    g�  �   �       �    ]�  �   �      �    ��  �   L      �    ;�  �   G      �    �C �          �    �%  �         �    4:  �   ]          5k  �   �       @    `T �   4           G�  �   K              �           #    �k  �   �      ,    �{  �   �      3     ` �           <    p$  �   Z      F    Yd  �   �       L    @0  �   A       S    2�  �   �       _    H�  �   2      f    ��  �   6      m    �.  �   �       u    �  �   2      |    �C �          �    C�  �   �       �    �(  �   �       �    i�  �   �       �    ��  �   �       �    � �   �       �    D�  �   O       �    � �   5      �    �  �         �    �0  �   i       �    ��  �   l      �    [ �   P       S    ��  �   �       �    �  �   5      �    b/  �   �       �    ��  �   z       �    j8  �   �      i     � �               ��  �   �           k�  �   Y           z�  �         %    �Y  �   9       4    6K  �   �      =    p �   �      1    � �   9       B    �C �          H       �          s
    �@ �           Q    HL �          W       �           ^    �C �          g     � �           m    z�  �   �       t    �4  �   9       ~    �1  �   g       �
     �   D       �	    t �   '       �    � �   >       �    � �   T       �    t�  �   V       �    ��  �   �       �    ?1  �   U       �    qi  �         �    � �   n       �    z�  �   }       �    �h  �   �       �    ڱ  �   �       �    � �   9       �    @D �          �    ��  �   S       	    �m  �   j      
	    �g  �   k       	    �<  �         t
    �@ �           !	    #�  �   W       (	    �R  �   H      3	    k�  �   �       :	    7�  �   �       A	    �g  �   �       M	    �H  �          X	    &a  �          c	    - �   X       m	    �-  �   �       t	    bJ  �   �       �    z�  �   D      �	    �  �   ]       �	     4 �          �	    @  �   D      �	    PL �          �	    K3  �   �      �	    �  �   �       �	    f�  �   �       
       �           �	    ��  �   9       �	     �   ;       �	    x�  �   b       �	    �C �          �	    <"  �   �      �	    �  �   K       �	    J �   *       �	    Ǖ  �   �       �	    ��  �   K       
    ��  �   �           � �   /       �
    D �          
    �)  �   r       
       �           
    �C �          �    ��  �   �       �    F �   a       '
    �]  �         �
    ��  �   S       0
    kw  �   +       �    ,  �   �      >
    �'  �   �       F
    ��  �   l       ?    *  �         P
    p�  �   �       y
    b �   9       W
    �z  �   I       ]
    9�  �   X       f
    �T  �   e      r
    �@ �           x
    s �   9       }
    ��  �   K       �    y�  �         �
    �o  �         �
    � �   Z       �
    ��  �   6      �
    � �   9       �
    
 �   �       �
    � �   2       F    ��  �   �       �
    �C �          �
    %O  �   i      �
    ��  �   �       �
    �&  �   �       �
    \Z  �   '          ��  �   �       
       �           �     D �          �
    }�  �   S       �
    9(  �   p       �
     0 �   @      �
    N   �                Ee  �   C          @ �   :           ��  �   u          d�  �   �       !    w�  �   ]       (    ��  �   �      4    D �          h     � �           =    F�  �   k       D    �  �   \      L    �  �   L       S    1�  �   Y       [    ��  �   �       �       �           e    &b  �   �       o    6�  �   7       t    D �          {    1�  �   �       �    ;Y  �   a       �    @�  �   U       '    +v  �         �    �Y  �   �       �    `L �          6    �q  �   �      �    �1  �   i       �    � �   ;       �    ��  �   3      �    `   �   �      �    �p  �   �       �    �  �   L       �       �           �    o�  �   U       �    2w  �   9       �    d2  �   �       �    Ð  �   �           z �   '       �       �               �5  �   ^           2�  �   �           c �   4       #    �  �   a       *    v�  �   �       0    � �   9       5    ��  �   +      ?    3�  �   D      L    O �   =       R    h�  �   �      [    ��  �   r       c    �0  �   U       o    ��  �   L       t    
c  �   O       lib/setup.asm HEADER_MAGIC HEADER_FLAGS header crt0.c explore.c .LC0 .LC1 file.c cfs.c .LC2 alloc_spin_lock pipe.c path.c gui.c font8x16.c window.c bmp.c font.c border.c editbox.c editbox_refresh mouse.c menubox.c obj.c objm foc message.c dialog.c button.c listbox.c file_data file_type file_unidade attr .LC3 .LC4 .LC5 .LC6 .LC7 .LC8 .LC9 .LC10 memcmp.c memcpy.c memset.c strcasecmp.c strcat.c strchr.c strcmp.c strcpy.c strcspn.c string.c strlen.c strncasecmp.c strncmp.c strncpy.c strpbrk.c strrchr.c strsep.c strspn.c strtok.c last.1481 strstr.c strdup.c memmove.c strcoll.c strerror.c ctype.c tolower.c toupper.c stdio.c fopen.c fclose.c fflush.c fputc.c fgetc.c fgets.c fputs.c fread.c fwrite.c remove.c rewind.c fseek.c feof.c ftell.c vfprintf.c vf vsprintf.c vsnprintf.c sn_buf putchar.c sscanf.c perror.c vfscanf.c character _buf.1638 fvalue _buf.1650 ungetc.c getchar.c freopen.c tmpnam.c _tmpnam rename.c itoa.c i2hex.c malloc.c calloc.c free.c realloc.c lldiv.c strtol.c atoi.c atol.c strtoul.c exit.c getenv.c qsort.c qscmp qses qsexc qstexc qs1 system.c strtod.c ftoa.c _precision atof.c strtof.c strtold.c abs.c ltoa.c utoa.c srand.c errno.c gmtime.c localtime.c strftime.c clock.c math.c pow.c sqrt.c atan.c acos.c asin.c floor.c ceil.c exp.c locale.c signal.c setjmp.c _GLOBAL_OFFSET_TABLE_ longjmp read_directory_blk menumotor drawstring strcpy log sqrt setjmp put clean_blk_enter strtok_r stdout vsprintf ungetc pwd_ptr argv strerror utoa_r __m_i memmove __tm __realloc_r atol __window_puts getenv ceil errno floor strtold _infinity loop qsort fgets file_update file_read_block m_file_list memcpy __window_clear BitMAP2 perror ltoa_r tolower system feof malloc remove fs_directory msg_read __window_putchar ldexp vsnprintf m_edit strtoul itoa __pipe__ stdgetc_r update_directory_entry _drawline fflush argc drawrect BitMAP eh_frame stdputc_r upath tell_r strncasecmp border button write_r strtol user rename flush_r strrchr update_editbox utoa calloc strtod fmouse rewind_r dialogbox atof update_objs seek_r strcat read_directory_entry debug_o fseek obj_focprocess __free_block_r open_dir ftoa stdin font8x16 __m_c _start obj_list __end strstr write_blk get_file_name atan2 signal strcoll strncmp write_sector draw_char_transparent pow strncpy put_pixel strcasecmp log10 _BLK_ realloc drawchar path_count open_file_r strtok remove_blk memcmp sscanf getfilename file_close pipe_write sigaction read_r file_write_block fread _ctype open_file addr search_blk_null strdup fopen sysgettmpnam localtime memset pwd main ftell srand init_process fclose getchar close_r __data ptr_mouse2 __free_r update_window getkeyw _vsputs_r strcmp color msg_init remove_file __bss atan fgetc drawchar_trans strtof strcspn asin ltoa setlocale stderr create_file strsep getkey __malloc_r fputc open_r A__ call_function getpathname strftime i2hex lldiv fwrite obj_process __window getmsg vfscanf rewind freopen msg_write pipe_read exit pipe_r register_obj __block_r atoi __heap_r ptr_obj assert_fn gmtime strspn ctr0 drawstring_trans strlen __code toupper wcl filename_cmp submenubox clock read_super_block abs strchr fputs acos strchrnul file_listbox frexp vfprintf strpbrk read_sector free setpath  .symtab .strtab .shstrtab .text .data .got .got.plt .data.rel.local .bss .eh_frame .comment                                                                                        �                                       !                �                                          '              @ �    @     p                              ,             p@ �   p@                                  5             �@ �   �@                                   E             �@ �   �@     @                             J              ` �    P      0                             T      0                �     *                                                   0�     �-      
   �                 	                      ح     |                                                   T�     ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ELF          >       �   @       ��         @ 8  @                   �      �                                      �      �   �        @                   P      ` �    ` �    0       0             Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��  ���_ cole _          �      �            � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           I��H�D �   L�H��C �   H�H�   �   L�H�  �   L�#H�  �   L�+�   �����H��H��H��H��L�������UH��AWSH��@��H�����I�      L�H�}�H�u�H�U�H�M�L�E�L�M�H���������H�H�U�H�H��     H�E�H�H�E�H�`     H�H�`     H�H� H��H��     H�H��     H�H��H�P     H�H�`     H�H�@H��H�H     H�H�E�H�h     H�H�E�H�@     H�H�E�H��     H�H��     H�H��H�X     H�I�߸    H��c������H���H�p     H�    H���������H�H� H��H�x     H�H���������H�H� H��H���������H�H� H�։�I��H���������H��ЉE�E��I��H�Z�������H��АH��@[A_]���UH��AWSH��0��H�����I�%     L�H�}�H���������H�4H��     H�<I��H���������H���H�E�H�}� u������rH�Eȋ@4�E�H�E�H�@8H�E؋U�H�M�H�Eؾ   H��I��H���������H���H�E�H��I��H�k�������H���H�E�H��I��H� �������H��и    H��0[A_]���UH��AWSH�� ��H�����I�?     L�H�8     �    H��jj j�A�/ A��  ��  �(   �   H���������H�<I��H�`�������H���H�� H�E�j�u�A�����A�    ��  ��  �    �    I��H�3������H���H��H�0     H�H�0     H�H��I��H��������H���H�u�H�E�jjA�(   A�    �    H�	�������H�H��I��H��������H���H��H�E�   H��������H�4H��I��H�|������H���H�E�   H��������H�4H��I��H�|������H���H�E�   H��������H�4H��I��H�|������H���H�E�   H�"�������H�4H��I��H�|������H���H�u�H�E�j jA�(   A�    �0   H�(�������H�H��I��H��������H���H��H�E�H��I��H��������H���H�E�H��I��H��������H���H�E�H��I��H���������H���H�0     H�H��I��H��������H���H���������H�H� �   H���rH�E�H��H�}�������H�������UH��AWSH�� ��H�����I�t     L�H�}�H�E�H�ƿ    I��H��������H��ЉE�E������   ��H��    H�G H�H�< H�>��H�8     ���u[H�E�H��     H�4H��I��H�J������H���H�8     �   H�0     H�H��H���������H����$H�0     H�H��H���������H������H�� [A_]���UH��H��0��H�����I�`     L�H�}�H�u��U܉M�L�E�H���������H�H� H�E��E�H9E�}?H�E��@��H9E�}0H�E�H�E��E�H�E�H��H�E�H�H��    H�E�HE؉������UH��SH��@��H�����I��     Lۉ}ԉuЉỦM�L�E�L�M�f�E�  H�E�H�@H�E�H�E��@�E�}�u�E�    �E�    �   f�E� H�E��@�EȉE��H�H� H�E�H�� f�E�H�E�� ���E��J�E�f#E�f��t5�UЋE��Hc��UԋE��H�H�}��M�U�I��H��H���������H���f�e�m��}� y��E�H�E��@9E��b�����H��@[]���UH��AWSH��0��H�����I��     Lۉ}܉u؉UԉM�D�E�L�M��E�    �X�E�    �CH�E�L��   �M�H�E��P�u؋E��Hc��}܋E��H�H��I��H���������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I�     Lۉ}܉u؉UԉM�D�E�L�M��E�    �p�E�    �[H�E�H��   �E��E�i��E��A��H�E��P�M؋E��Hc��M܋E��H�I��D��H��I��H���������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I�<     Lۉ}܉u؉UԉM�D�E�L�M��}� �[  �}� �Q  �E�    �>H�E�L��   �M�H�E��P�E�Hc��}܋E��H�H��I��H���������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E����Hc��}܋E��H�H��I��H���������H��ЃE��E�;E�|��E�    �AH�E�H��   �M�H�E��P�u؋E��Hc��E�H�I��H��I��H���������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E��Hc��}܋E����H�H��I��H���������H��ЃE��E�;E�|���H��0[A_]���UH��AWSH��@��H�����I��     Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}��  �E�    ��   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��   �E�f#E�f��tDH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H���������H����BH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H���������H���f�e�m��}� �[����E�H�E��@9E��	�����H��@[A_]���UH��SH��8��H�����I�*     L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H�_�������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I�l     Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}���   �E�    �   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��W�E�f#E�f��tBH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H���������H���f�e�m��}� y��E�H�E��@9E��T�����H��@[A_]���UH��SH��8��H�����I�O     L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H���������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I��     L�H�}ȉuĉU��M�D�E�D�M�H���������H�H� H�E�H�E�H   � �? �    H��I��H��s������H����E�    �U�H�E��P4�UH�E��P8�UH�E��P<H�E��@H   H�E��@L   H�E��P<H�E��PP�UH�E��PTH���������H�H��H�E�H�PXH�E��@D    H�E��PDH�E��P@�U�H�E��P�U�H�E��P�U�H�E��P �U�H�E��P�U H�E��P`�} u�E�   H�E��@�P�H�E��P(H�E��P�E�)ЍP�H�E��P$H�E��@0   �E����H�E��P,H�E��@��H�E��@��H�E�I���Ѻ    �    I��H� ������H���H�E��@4��H�E��@����H�E�I��A�ȹ   �   �   H�?�������H��Ѓ}� u:H�E��@����H�E�I��A���� �   �   �   H�?�������H����8H�E��@����H�E�I��A���� �   �   �   H�?�������H��Ѓ}� t}H�E��@����H�U��E�I��A���� ����   �   H�?�������H���H�E��@4��H�E��@���ƋE��H�U�I��A�ȹ   ��ƿ   H�?�������H���H�E��@8A��H�E��@$��H�E��@(��H�E��@,��H�E��@0��H�E�I��H�?�������H���H�E�H��I��H�
y������H������E�H�E�H�pHH�E��@��E܉������)Љ�H�E�H���u�I��A���� ������   ��H��H���������H���H��H�E��@����H�E�I��A�    �   �   �   H���������H���H�E�H�PHH�E��@��H���u�I��A���� ������   �ƿX   H���������H���H��H�E�H�PHH�E��@��(H���u�I��A���� ������   �ƿ-   H���������H���H��H�E�H�e�[A_]���UH��AWSH��0��H�����I�     L�H�}�H�u�H�E��P0H�E��@Ѓ�P�E�H�E��P,H�E��@Ѓ��E��E�P   �E�   �E�    �E���� H�E�H��I��H�
y������H��ЉE�H�E�L�@H�M؋U܋E���������p��E�<�E��������ƋE���)ƋE��H�E�H���u�M��A�ȉщ�H��H���������H���H���H�e�[A_]���UH��H����H�����I�	     L�H�}��   H�E�H���r�����UH��H����H�����I��
     L�H�}������UH��H����H�����I��
     L�H�}�H�U��BD    H�U��JDH�U��J@H�U��R8A��H�U��R$��H�U��R(A��H�U��R,��H�U��R0��H�U�I��D��I�?�������J��А����UH��SH��(��L�����I�
     Mډ�f�E�H���������I�H� H�E�H���������I�H��H�E�H�PXH�E�@(�P�H�E�@H���к    ��E�H�E�@$�P�H�E�@L���к    ��E�H�E�P<H�E�PPH�E�PD�E�9�rH�E��@D    H�E�@@�PH�E�P@H�E�P@�E�9�r9H�E��@D    H�E�PDH�E�P@H�E�H��H�O�������I����E��  f�}���   H�E�@D����   H�E�@D�P�H�E�PDH�E�H�xHH�E�pTH�E�@PH�U�J,H�U�RLA��H�U�R@A��ʃ���H�U�J0H�U�RHA��H�U�RDA��ʃ�A��H���u�I��A������D�޿    H�_�������I���H����   f�}�	uH�E�@D�PH�E�PD��   f�}�
u!H�E��@D    H�E�@@�PH�E�P@�   f�}���   H�E�H�xHH�E�pTH�E�PPH�E�H,H�E�@LA��H�E�@@A��ȃ���H�E�H0H�E�@HA��H�E�@DA��ȃ�A���E�H���u�I��A���щ�D�މ�H�_�������I���H��H�E�@D�PH�E�PD�E�H�]�����UH��H����H�����I�R     L؉}�H���������H�H� H�E��U�H�E��P<�����UH��SH��(��H�����I�     L�H�}�H�}� t=H�E�H�E��&H�E�H�PH�U�� f�����H���������H���H�E�� ��u���H��([]���UH��AWSH��P��H�����I��     L�H�}��u��U��M�L�E�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H���������H�<I�߸    H�f�������H��Ҹ�����6  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H���������H�<I�߸    H�f�������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H���������H�<I�߸    H�f�������H��Ҹ   ��   �E�    �   �E�    �   �}� tNH�E�H��   H�E��P�M��E���E��Hc��M��E���E��H��M�I��H��I��H���������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H���������H��ЃE��}� �U����E��}� �;����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��P��H�����I��     L�H�}��u��U��M�D�E�L�M�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H���������H�<I�߸    H�f�������H��Ҹ�����3  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H���������H�<I�߸    H�f�������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H���������H�<I�߸    H�f�������H��Ҹ   ��   �E�    �   �E�    �   �}� tKH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H���������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H���������H��ЃE��}� �X����E��}� �>����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��0��H�����I��      Lۉ}܉u؉U�H�M��E�    �   �E�    �t�U�������E��H���������H�Hڋ��E�}� tBH�E�H��   H�EȋP�MԋE��Hc��M؋E��H��M�I��H��I��H���������H��ЃE��}�~��E��}��o�����H��0[A_]���UH��AWSH��@��H�����I���      Lۉ}̉uȉUĉM�L�E��E���� �E�``` �E���� �EĉE��ẺE܋E��E؋EȉEԋE؍P��E��xH�M��E�I��A�    �   ��I��H���������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H���������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H���������H��ЋEԍP��E܍pH�M��E�I��A�    �Ѻ   ��I��H���������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H���������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H���������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H���������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H���������H��ЋEԍP��E܍p�M��E�ȃ�H�M�I��A�    �Ѻ   ��I��H���������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H���������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H���������H��ЋE؍P��M܋E�ȍp��E���H�M�I��A�    �   ��I��H���������H��АH��@[A_]���UH��AWSH��0��H�����I���      Lۉ}܉u؉UԉM�D�E�D�M�H�} u
�    ��  �H   I��H��������H���H�E�H�}� u
�    ��  H�E�H   �    H��I��H��s������H���H�UH�E�H�P@H�E�U�PH�E�P0�E��H�E�PH�E�P,�E��H�E�PH�E��    H�E�P(�E�9�wH�E�P(H�E�P�
�U�H�E�PH�E�P$�E�9�wH�E�P$H�E�P�
�U�H�E�P�U�H�E�P�U�H�E�P H�E��@0    H�E�@0��I��H��������H���H��H�E�H�P8H�E�H�@8H��t.H�E�@0H�U�H�R8H�щ¾    H��I��H��s������H���H�E�@ ��H�E�@��H�E�@��H�E�@��H�E�@L�MA����I��H�?�������H���H�E�@��H�E�@��H�E�@��H�E�@L�MA�������I��H���������H���H�E�H��0[A_]���UH��AWSH�� ��H�����I�z�      L�H�}�H�E�H�@@H�E�H�E؋@ A��H�E؋@��H�E؋@��H�E؋@��H�E؋@��H�E�I��I��H�?�������H���H�E�H��H��������H��АH�� [A_]���UH��AWSH�� ��H�����I���      L�H�}�H�}� u
������z  I�߸    H��0������H��҉E�}���   I�߸    H��0������H��҉E�}�[��   I�߸    H��0������H��҉E�}�Ct�}�Dt'�GH�E؋P,H�E؋@49�s1H�E؋@,�PH�E؉P,�H�E؋@,��tH�E؋@,�P�H�E؉P,����H�E�H��H��������H��и    �  H�E�H�P8H�E؋@,��H�H�E��}� �C  H�E؋P,H�E؋@09��-  H�E��@    �}���   H�E؋@4��tkH�E؋@,��t`H�m�H�E؋P4H�E؋@,)�H�E�H�HH�E�H��H��I��H�ր������H���H�E؋@,�P�H�E؉P,H�E؋@4�P�H�E؉P4�   H�E��@   �~H�E؋P,H�E؋@49�t4H�E؋P4H�E؋@,)�H�E�H�HH�E�H��H��I��H�ր������H��ЋE��H�E��H�E؋@,�PH�E؉P,H�E؋@4�PH�E؉P4H�E��@   H�E�H��H��������H���H�E؋@����u*H�E�H��H��������H���H�E؋@����H�E؉P�    H�� [A_]���UH��AWSH��@��H�����I��      L�H�}�H�E�H�@@H�E�H�E�H�@8H�E��E�    f�E�  H�E��@��uH�E��@    �  �E�    �  �E�    �E�    ��   �}� ueH�E��P4�E�9�vH�E�H�PH�U�� f�f�E��f�E�  f�}�
uf�E�  �E�   H�E��P,�E�9�u�U�H�E��P$�U�H�E��P(�E�f�}� teH�E�H�xHH�E��p H�E��PH�E��H�E��A��H�E��H�E��A���E�H���u�I��A����D��D�։�I��H�_�������H���H���E�H�E��P�E�9������E�H�E��P�E�9������H�E�H�xHH�E��p H�E��@H�U��JH�U��R(�A��H�U��JH�U��R$�A��H���u�I��A����D��D�ֿ_   I��H���������H���H��H�e�[A_]���UH��AWSH��@��H�����I��      L�H�}�H�E��@ �E�H�E��@�E�H�E��@�E�H�E��@�E�H���������H�H� � �E�H���������H�H� �@�E�H���������H�H� �@�E̋EЃ����X  �E�;E�~Q�E���9E�~F�U�E��9E�}9�E��P�E��9E�})�E�+E��E�+E�։�I��H�I������H�����   �E�;E���   �E�;E���   �U�E��9E���   �U��E��9E���   H���������H�H� � ��H�E��@ )ЉE�H���������H�H� �@��H�E��@)ЉE��aH���������H�H� � +EȉE�H���������H�H� �@+EĉE�}� y�E�    �}� y�E�    �U�H�E��P �U�H�E��PH���������H�H� �@����u�I�߸    H�3������H��ҐH��@[A_]���UH��AWSH��@��H�����I���      L�H�}�H�u�H�UȉM�D�E�D�M��P  I��H��������H���H�E�H�E�P  �    H��I��H��s������H���H�E�H��I��H�
y������H��ЉE�}�~�E�   �U�H�E�H�H0H�E�H��H��I��H�%s������H���H�E��    H�E��U�P�U�H�E��P�E�����H�E��P�U�H�E��P�UH�E��PH�U�H�E�H�P(H�E�H�PHH�E��@����H�E��@����H�E�H��0H���u�I��A���� �    ��H��I��H���������H���H��H�E�H�U�H��H�e�[A_]���UH��AWSH��0��H�����I�u�      L�H�}�H�uЉU�H�E؋@$��H��H��H�H��H�PPH�E�H�H��H�E�H�E؋@$�HH�U؉J$H�U؉�H��H��H�H��H�H�PP�ẺH�E�H��I��H�
y������H��ЉE�}�~�E�   �U�H�M�H�E�H��H��I��H�%s������H��и    H��0[A_]���UH��AWSH��P��H�����I���      L�H�}��E�    �E�����H�E�H�@(H�E�H�E�H�PHH�E��@����H�E��@����H�E�H��0H���u�I��A���� �  � ��H��I��H���������H���H��H�E�H�PHH�E��@����H�E��@��H���u�I��A���� �  � ���H���������H�<I��H���������H���H��H�E؋P0H�E��@ЉE�H�E؋@,�E��E�d   �E�   �EĀ�� �E�    �H���������H�H� �@����u�H�E��@$���A  H�E��P$�E���A��H�}؋MċŰuЋE�I��A��D�щ�I��H�?�������H����E�    �  H���������H�H� � ��H�E؋@ )ЉE�H���������H�H� �@��H�E؋@)ЉE�H���������H�H� �@�E�E�Hc�H��H��H�H��H�PPH�E�H�H��H�E��E�;E���   �E��E��E�Ѓ�9E���   �UԋE��9E�}�E��E��E�E��9E�}gH�E�H�xH�MċE��E��E�ЍP�EԍpH�E�H���u�I��A�ȹ����H��I��H���������H���H���E��E�m��E����tZ�nH�E�H�xH�MċE��E��E�ЍP�EԍpH�E�H���u�I��A�ȹ    H��I��H���������H���H���E������E�H�E��P$�E�9��[����E�����A����}��t5H�M��E�Hc�H��H��H�H��H�H��P� ��I��H�j������H����E�   �H���������H�H� �@����u�H�E�H�PHH�E��@����H�E��@����H�E�H��0H���u�I��A���� �    ��H��I��H���������H���H���E�H�e�[A_]���UH��AWSH����H�����I�q�      L�H�}�H�P       H�    H�X       H�    I�߸    H��������H���H�`       �    H�}� t'H�E� ��H�`       �H�X       H�E�H��    H��[A_]���UH��AWH����H�����I���      L�H�`       �����   ����   ��t
��tA�   H�X       H�H����   H�X       H�H��I��H�������H����yH�X       H�H��tbH���������H�<I�׸    H�f�������H����?H�X       H�H��t+H�X       H�H��I��H�0'������H����������    H��A_]���UH��AWSH��@��H�����I���      Lۉ}��u�H���������H�H� H��t�}� x�}� y&�H���������H�H� �@����u������#  H�E�    H�E�    �E�    �E�    �E�    �E�    �   H�P     �E�H�H�H��H�E�H�E�H��� �E�H�E�H��� �E�H�E�H��� �E�H�E�H��� �EċEԉE܋E�;E�~"�E�;E�~�UЋE��9E�}�ŰE��9E�|&�E��E�Hc�H���������H�H� H9��^������E�Hc�H���������H�H� H9�u&�H���������H�H� �@����u������  H�E� ���V  ����  ����  ���n  ��t����   �[  H�P     �E�H�H�H��H��H�P       H�H�P       H�H�@(H�E�H�P       H��@��I��H�j������H���H�P       H�H��I��H�c������H��ЉE���  H�P     �E�H�H�H��H��H�X       H�H�X       H�H�@@H�E�H�X       H��@��I��H�j������H����E�    H�`       �   �H���������H�H� �@����u��]  H�P     �E�H�H�H��H��H�X       H�H�X       H�H�@@H�E�H�X       H��@��I��H�j������H����E�    H�`       �   �H���������H�H� �@����u���   H�P     �E�H�H�H��H��H�X       H�H�X       H�H�@@H�E�H�X       H��@��I��H�j������H����E�    H�`       �   �H���������H�H� �@����u��*�H���������H�H� �@����u��E�    ������I�}� t>��H�E�� ��u�H�E�� �PH�E��H�E�H��H��������H���H�E��     �    H��@[A_]���UH��AWSH����H�����I��      L�H�}�H���������H�H� H��u*�   �    H�P     H�<I��H��s������H���H���������H�H� H=�   ~�    �LH���������H�H� H�HH���������H�H�
H�U�H�P     H�H��H���������H�H� H��[A_]���UH��AWSH�� ��H�����I�'�      L�H�}�H�E�    H�E؋@8A��H�E؋@$��H�E؋@(��H�E؋@,��H�E؋@0��H�E�I��I��H�?�������H����E�    �   H�P     �E�H�H�H��H�E�H�E�� ��tWH�E�� ��uOH�P     �E�H�H�H��H��H�X       H�H�X       H�H��I��H�w������H��������E��E�Hc�H���������H�H� H9��\�����H�� [A_]���UH��AWSH�� ��H�����I���      Lۉ}�H�u�H�E�H��I��H��
������H��и    H�.������H��҉E�E�H�� [A_]���UH��H����H�����I���      L؉}�H�P     ���	v5H�P     �D    H�P     �    H�P     �D    H�P     ��JH�P     �0�M�H�P     ��H�0�L�H�P     �T�JH�P     �L�����UH��H����H�����I���      L�H�P     �T��u
�    �   H�P     �T��	vH�P     �D    H�P     �LH�P     ��HT��U�H�P     �T�JH�P     �L0H�P     ��H��D�    �E�����UH����H�����I��      L�H�P     �D    H�P     �    H�P     �D    �]���UH��AWSH��0��H�����I���      L�H�}�H�u�H�E�H�E�H�Eȋ@��-�   �E�H�Eȋ@���2�E��E�,  �E�d   �EԍH��E؍P��E܍p�E���H�}�I��A�  ��I��H�?�������H��ЋEԍH��E؍P��E܍p�E���H�}�I��A�������I��H���������H���H�}ȋMԋU؋u܋E�I��A�������I��H���������H���H�E�H�HH�E܍P�E���
H���u�I��A�    �������H���������H�<I��H���������H���H���E��E��m��m�J�EԍH��E؍P��E܍p�E���H�}�I��A�������I��H�?�������H��ЋEԍH��E؍P��E܍p�E���H�}�I��A�������I��H���������H���H�}ȋMԋU؋u܋E�I��A�������I��H���������H����E�    I�߸    H��0������H���f�E�f�}�
��   f�}� tl�}� ~ff�}�u_�m�f�E�  H�E�H�xH�E܍P�E��H�E����4�E�H���u�I��A������    ��I��H�_�������H���H��H�m��of�}� �\���H�E�H�xH�E܍P�E��H�E����4�E�H���u�I��A������    ��I��H�_�������H���H���E�H�E�H�PH�U��U҈������H�E��  ��H�Eȋ ��u�H�Eȋ �PH�EȉH�E�H��I��H��������H���H�E��     �    H�e�[A_]���UH��AWSH��0��H�����I�;�      L�H�}��E���� �E�``` �E���� H�Eȋ@0��(�E�H�Eȋ@,��d�E��E�d   �E�2   �E؍P��E��xH�MȋE�I��A�    �   ��I��H���������H��ЋE؍P��E܍p�E���H�}ȋM�I��A�ȹ   ��I��H���������H��ЋE؍P��E܍p�E���H�}ȋM�I��A�ȹ   ��I��H���������H��ЋEԍP��E܍pH�MȋE�I��A�    �Ѻ   ��I��H���������H��ЋEԍP��E܍p�E���H�}ȋM�I��A�ȉѺ   ��I��H���������H��ЋEԍP��E܍p�E���H�}ȋM�I��A�ȉѺ   ��I��H���������H��ЋEԍP��E܍p�M��E�ȃ�H�}ȋM�I��A�ȉѺ   ��I��H���������H��ЋEԍP��E܍p�M��E�ȃ�H�}ȋM�I��A�ȉѺ   ��I��H���������H��ЋEԍP��E܍p�M��E�ȃ�H�M�I��A�    �Ѻ   ��I��H���������H��ЋE؍P��M܋E�ȍp��E���H�}ȋM�I��A�ȹ   ��I��H���������H��ЋE؍P��M܋E�ȍp��E���H�}ȋM�I��A�ȹ   ��I��H���������H��ЋE؍P��M܋E�ȍp��E���H�M�I��A�    �   ��I��H���������H��АH��0[A_]���UH��AWSH��0��H�����I��      Lۉ}܉u؉UԉM�D�E�D�M�H�} u
�    ��  �H   I��H��������H���H�E�H�}� u
�    ��  H�E�H   �    H��I��H��s������H���H�UH�E�H�P@H�E�U�PH�E�P0�E��H�E�PH�E�P,�E��H�E�PH�E��    H�E�P(�E�9�wH�E�P(H�E�P�
�U�H�E�PH�E�P$�E�9�wH�E�P$H�E�P�
�U�H�E�P�U�H�E�P�U�H�E�P H�E��@0    H�E�@0��I��H��������H���H��H�E�H�P8H�E�H�@8H��t.H�E�@0H�U�H�R8H�щ¾    H��I��H��s������H���H�E�@ ��H�E�@��H�E�@��H�E�@��H�E�@L�MA����I��H�?�������H���H�E�@��H�E�@��H�E�@��H�E�@L�MA�������I��H���������H���H�E�H��0[A_]���UH��AWSH��0��H�����I���      L�H�}�H�}� u
������,  I�߸    H��0������H��҉E�}���   I�߸    H��0������H��҉E�}�[uqI�߸    H��0������H��҉E�}�At�}�Bt �2H�Eȋ@,��t&H�Eȋ@,�P�H�EȉP,�H�Eȋ@,�PH�EȉP,��H�E�H��H��(������H��и    �pH�E�H��I��H���������H���H�E�H�EȋP(H�E�� 9�s=H�E�� ��H�EȉP(H�Eȋ@(��:vH�E��@(    H�E�H��H��(������H��и    H��0[A_]���UH��AWSH��@��H�����I�P�      L�H�}�H�E�H�@@H�E�H�E�H�@8H�E�H�E�@   H��H��������H�<I��H��T������H��ЉE��E�    H�E��@���E���H�EЋ ��u�H�EЋ �PH�EЉ�E�    �!  H�E��@�E�H�E��@ �E�H�E��P,�E�9�u�E�i� �E�����H�E��@��A��H�E��@�U���Ѓ���H�E��@����H�UЋE�I��A���   D��I��H�?�������H��ЋE�;E���  H�E�H��H��+������H���H�E�H�xH�u؋U�H�E��@�M���ȃ�A��H�E��H�E�ȃ�A��H�E�H���u�I��A����D��D��H��I��H���������H���H��H�E��@��E�ЉE�H�E�H�xH�u؋E�H�U��R�M���ʃ�A��H�U��J�U�ʃ�A��H���u�I��A����D��D��H�p       H�<I��H���������H���H��H�E��@���E�ЉE�H�E�H�xH�u؋E�H�U��R�M���ʃ�A��H�U��J�U�ʃ�A��H���u�I��A����D��D��H��       H�<I��H���������H���H���E�    H�m考E��E�;E������H�E��     �H�e�[A_]���UH��AWSH��@��H�����I�`�      L�H�}�H�E��@b���� ����  H��������H�H��������H�4H��       H�<I�߸    H���������H���H�E��@o��H��x�H*��H��H���H	��H*��X��E�H�(���������E��E�    H�E��@o=���?v�E�   H�0���������E��)H�E��@o=�� v�E�   H�8���������E��E��^E��E�H�E�fHn�H��������H�4H�p       H�<I�߸   H���������H���H�p       H�<I��H�
y������H��ЉE̋ẺE��H�p       �E�H�H�� �E��}�~�H�        �E�H�H�H��H�w       H�H��������H�4H��I�߸    H���������H����   H�#�������H�H��������H�4H��       H�<I�߸    H���������H���H�#�������H�H��������H�4H�p       H�<I�߸    H���������H��ѐH��@[A_]���UH��AWSH����H�����I���      Lۉ}�H�u�H�E�� ��H�E��@9�sH�E��P#H�E��@9�r"H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@��u)H���������H�H��E�H�։�H�$.������H���H�E�H�PH�E��@#��H�H�E�H�PH�E�H�@�U�H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  H�E��@��u0H���������H�H� H��t�E�����I��H���������H��ЋE�H��[A_]���UH��H����H�����I�v�      L�H�}��E�    H�E�@��u]H�E�@'�PH�E�P'��H�E�P#H�E�@'9�r�H�E�H�PH�E�@'��H��H�H�E�H�PH�E�H�@� ���E��   H�E�@��tH�E�@��uiH�E�@#��u������ZH�E�P'H�E�@#9�r������AH�E�H�PH�E�@'��H�H�E�H�PH�E�H�@� ���E�H�E�@'�PH�E�P'�E�����UH��H����H�����I�X�      L�H���������H�H� H�E��E�    H�E��@��uWH�E��P#H�E��@'9�w�    �AH�E�H�PH�E��@'��H�H�E�H�PH�E�H�@� ���E�H�E��@'�PH�E��P'�E�����UH��H����H�����I���      L�H���������H�H� H�E��E�    H�E��@��uXH�E��@'�PH�E��P'��H�E��P#H�E��@'9�r�H�E�H�PH�E��@'��H��H�H�E�H�PH�E�H�@� ���E��E�����UH��AWH��(��H�����I��      L�H�}�H�u�H�U����u�    �(H�M�H�U�H��H��I��H��I������H���H�E�H�E�H��(A_]���UH��AWSH�� ��H�����I���      L�H�}�H�}� u
������   H�}� tH�E؋@����tH�E��@"<t������zH�E؋@%�   ��u�    �cH�E؋@#H�U؋J�    ��E�H�E؋@��@��u�U�H�E؉�H��I��H�T������H���H�E�H��I��H�Q������H��ЉE�E�H�� [A_]���UH��AWSH����H�����I���      L�H�}�H�}� u������0H�E�H��H�]2������H���H�E�H��I��H�BR������H���H��[A_]���UH��AWSH�� ��H�����I�;�      Lۉ}�H�u�H�}� u
�������  H�EЋ@��u
�    �  H�EЋ@��tH�EЋ@��tH�EЋ@��u!H�UЋE�H�։�H�$.������H����y  H�EЋ@����unH�EЋP#H�EЋ�+  9�wYH�EЋ�+  ��tKH�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��E�U�H�EЉ�H��I��H�BS������H����H�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U܈H�E�� ��H�EЋ@��9�r3H�EЋ@����H�EЉPH�E�f�   H�E�H��H�]2������H���H�EЋ@#�PH�EЉP#H�EЋP#H�EЋ�+  9�vH�EЋ�+  �PH�EЉ�+  H�EЋ@���H�EЉP�    H�� [A_]���UH��AWH��(��H�����I� �      L�H�}�H�}� u
������  H�E؋@��u
�    �v  H�E؋@��tH�E؋@��tH�E؋@��u"H�E�H��H�~/������H��ЉE�E��0  H�E؋P#H�E؋�+  9�r
������  H�E؋@����ulH�E؋P#H�E؋�+  9�wWH�E؋�+  ��tIH�E؋@����H�E؉PH�E؋@#H�U؋r�    ���E�U�H�E؉�H��I��H�BS������H���H�E؋@#H�U؋J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@� ���E�H�E�� ��H�E؋@��9�rH�E؋@����H�E؉PH�E�f�   H�E؋@#�PH�E؉P#�E�H��(A_]���UH��SH��H��H�����I�R�      L�H�}ȉuĉU�H�M�H�}� u�    �y�E�    H�E�H�E��E�    �FH�E�H��H��5������H��ЉE؃}��u�E�    �u��4H�E�H�PH�U��U؈�E��E��E��E��E�9�w��E�    �u�H��H[]���UH��SH��H��H�����I���      L�H�}ȉuĉU�H�M�H�}� u�    �l�E�    H�E�H�E��E�    �9H�E�H�PH�U�� ���E�H�U��E�H�։�H��3������H��ЃE��E��E��E��E�9�w��E�    �u�H��H[]���UH��H����H�����I���      L�H�}�H�u��U�}�tZ�}�|�}� t�}�t�nH�E���H�E��P#H�E���H�E��P'�RH�E��@#H�U��H�E��P#H�E��@'H�U��H�E��P'�(H�E���+  H�U�)Љ�H�E��P#H�E��P#H�E��P'�H�E��@#H�U��J�    ��Љ�H�E�f��    ����UH��H����H�����I� �      L�H�}�H�}� u�    �	H�E��@#������UH��H����H�����I���      L�H�}�H�}� t7H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@����H�E��P������UH��H��(��H�����I�V�      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H��(��H�����I��      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H����H�����I���      L�H�}��E�_   �(�E�Hc�H�E�H�� < u�E�Hc�H�E�H��  �m��}� y����    ����UH��H����H�����I�C�      L�H�}�H�E�H�E�H�E�H�E��H�E�� </uH�E�H��H�E�H�E�H�E�� ��u�H�E�����UH��H��0  ��H�����I���      L�H������H������H������H�E�H������H�E�H������H�E��E�    �?H�E�� ��u�E�Hc�H�E�H��  �H�E�H�PH�U��U�Hc�H�U�H�� ��E��}�_~��E�    �-H�E�H�PH�U��H�E�H�PH�U�� 8�t�   ��E��}�_~͸    ����UH��SH�� ��H�����I���      L�H�}�H�u�H�E؋PH�E؋@ЉE�E�H�U����H��     H�H�¾   H��:������H��ЉE�}� t
�������   �E�    ��   �E�%�  ��H��     ��H؋���uf�E�%�  ��H��     ��H��������E�H�U����H��     H�H�¾   H��:������H��ЉE�}� t������r�E��m�E�%�  =�  uE�E��E�H�U����H��     H�H�¾   H��:������H��ЉE�}� t�������E�H�E؋@$9E����������H�� []���UH��H����H�����I�k�      L؉}��u�H�U�H�M�    ����UH��AWSH��0��H�����I�/�      Lۉ}�H�u�H�U�H�EȋPH�Eȋ@ЉE�H�Eȋ@ �E܉E�ЉE�   �    H��     H�<I��H��s������H����E�    �B�U�E�Љ�H�EЋ ��H��     H��   H��:������H��ЉE��}� u�E�H�EȋP �E�9�w���H��0[A_]���UH��H����H�����I�I�      L�H�}�H�u�H�U��R��H�U����H�U�H��H��   I��:������J� ������UH��AWSH��`��H�����I��      L�H�}�H�u�H�U�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H��������H���H�E�H�E�H�E�H�E�H��I��H�<q������H��ЉE�H�E��@,�E��9  H�E�H�E��H�E�� </uH�E��  H�E��H�E�H�E�� ��u׋U�H�E��@ H�M��	��H�M���H��:������H��ЉE؃}� t#H�E�H��I��H���������H��и    ��   �E�    �f�E���Hc�H�E�H�H�E�H�E��@a��t5H�E��@b����@��t#H�E�H�U�H��H��H�<������H��ЉE���E������}� t�E��}�?~����}� u+�}�?%H�EЋ@k�E�H�E��@ �E؉E�ЉE�m��	�E�    �
�}� �����H�E�H��I��H���������H��ЋE�H��`[A_]���UH��AWSH��P��H�����I�ӽ      L�H�}�H�u�H�U��M�L�E�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H��������H���H�E�H�Eغ    �    H��I��H��s������H��ЋU�H�E��@ H�M��	��H�M؉�H��:������H��ЉE�}� t#H�E�H��I��H���������H��и������   �E�    �T�E���Hc�H�E�H�H�E�H�E��@a��t#H�E�H�U�H��H��H�<������H��ЉE���E������}� t�E��}�?~����}� u:�}�?4�E���Hc�H�E�H�H�EȺ�   H��H��I��H�%s������H�����E�����H�E�H��I��H���������H��ЋE�H��P[A_]���UH��AWSH��P��H�����I�	�      L�H�}�H�u�H�U�H�E���C  ��u
������	  H�E���C  ��@v/H�@�������H�<I�߸    H�f�������H��Ҹ������  H�E��PH�E��@ЉE�H�E���?  H�E��@ �ЋE�ЉE�    I��H��������H���H�E�H�Eغ    �    H��I��H��s������H��ЋU�H�E��@ H�M��	��H�M؉�H��:������H��ЉEԃ}� t!H�E�H��I��H���������H��ЋE��  H�E���C  ��H��H��H�E�H�H�E�H�EȺ`   �    H��I��H��s������H���H�E�H��+H��H��;������H���H��H�E�H��H��I��H�.v������H����E�    �"H�UȋE�H����uH�UȋE�H�� �E��}�_~�H�E��@` H�E���+  H�EȉPo�U�H�E��@ H�M��	��H�M؉�H��:������H��ЉE�H�E�H��I��H���������H��ЋE�H��P[A_]���UH��AWSH��`��H�����I���      L�H�}�H�u�H�U��S  I��H��������H���H�E�H�EкS  �    H��I��H��s������H���H�E��PH�E��@ ��H�EЉP�    I��H��������H���H�U�H�BH�E��PoH�EЉ�+  H�E��PH�EЉ�/  H�E��P H�EЉ�3  H�E��H�EЉ�G  �    I��H��������H���H�U�H��K  H�E�H��K  �    �    H��I��H��s������H���H�E��@k�E�    I��H��������H���H�E��E������E�    �E�    ��  �   I��H��������H���H�U�H��K  �M�Hc�H��H�H�H�E�H��K  �U�Hc�H��H�H� H�E�H�E��   �    H��I��H��s������H����E�    �<  H�E��@ �E��H�E��@�H�E��P�E�H�H�4�    H�E�H�ʉH�EЋ�;  �PH�EЉ�;  �E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E�;E�ts�E�H�U����H�U�H��H�¾   H��:������H��ЉE��}� t:H�E�H��I��H���������H���H�E�H��H�BR������H��и    �   �E��E�H�E��@�����E�    ��U�E�H��    H�E�HЋ �E�}��u	�E�������E��}��  ������}��t�E��}��  � �����H�E�H��I��H���������H���H�E�H��`[A_]���UH��AWSH��p  ��H�����I�*�      L�H������H�������   I��H��������H���H�E�H�E�H�E�H�E�H   H�E�H������H�E�H��H��I��H��n������H���H�U�H�E�H��H��I��H��q������H��п�   I��H��������H���H��     H�H��     H���   �    H��I��H��s������H��п   I��H��������H���H�E�H�EȺ   �    H��I��H��s������H���H�E�H�E�H�E��   �    H��I��H��s������H����E�    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ ���    Hǅ���    Hǅ���    Hǅ���    Hǅ ���    Hǅ(���    Hǅ0���    Hǅ8���    Hǅ@���    HǅH���    HǅP���    HǅX���    Hǅ`���    Hǅh���    Hǅp���    Hǅx���    H�E�    H�E�    H������H������H��H��I��H�.v������H���������<wt������<au�E�   H�E��@   H�E��     H�U�H�E�H��H��H��?������H��ЉE�}� t_H��     H�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��и    �  H�E�H�U�H�M�H�E�H��H��H�	@������H��ЉE��}� u_H��     H�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��и    �  H�EȋU��P,H��     H�H�M�H�U�H�u�I�ȹ    H��H�B������H��ЉE�}����   �}� tqH��     H�H������H�U�H�u�A�    H��H��X������H���H��     H�H������H�U�H�u�I�ȹ    H��H�B������H��ЉE�}� ��   H��     H�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��и    ��  �}� t_H�E�H��I��H���������H���H��     H�H��I��H���������H���H�E�H��I��H���������H��и    �r  H��     H�H�U�H�M�H��H��H�EF������H���H�E�H�}� ��   H��     H�H��H�E�H��+�`   H��H��I��H�%s������H���H�E�H��+H��H�H;������H���������<wt������<+t������<au
H�E��@"�H�E��@"H�E��@   H�EȋP,H�E���?  H��     H��PsH�E���C  ������<auH��     H��PoH�E��P#H�E�H��I��H���������H���H��     H�H��I��H���������H���H�E�H��I��H���������H���H�E�H��p  [A_]���UH��AWSH��@��H�����I��      L�H�}��   I��H��������H���H�E�H�E�   �    H��I��H��s������H���H�E�H�E�H�E�   �    H��I��H��s������H���H�E��@   H�E��     H�U�H�E�H��H��H��?������H��ЉE܃}� t H�E�H��I��H���������H��и�����AH�U�H�M�H�E�H��H��H��C������H��ЉE�H�E�H��I��H���������H��ЋE�H��@[A_]���UH��AWSH�� ��H�����I���      L�H�}�H�E�H�@H��I��H���������H����E�    �TH�E�H��K  �U�Hc�H��H�H� H��t?H�E�H��K  �U�Hc�H��H�H� H��I��H���������H��ЃE��}��  ~���H�E�H��K  H��I��H���������H���H�E�H��I��H���������H���H�E�    �    H�� [A_]���UH��H�� ��L�����I���      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H��:������I� ������UH��H�� ��L�����I�ޫ      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H��:������I� ������UH��AWSH��   ��H�����I��      L�H��x���H��p�����l����   I��H��������H���H�E�H�E�H�E�H�E�H   H�E�H��x���H�E�H��H��I��H��n������H���H�U�H�E�H��H��I��H��q������H��п   I��H��������H���H�E�H�EȺ   �    H��I��H��s������H���H�E�H�E�H�E��   �    H��I��H��s������H���H�E��@   H�E��     H�U�H�E�H��H��H��?������H��ЉE��}� t_H��     H�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��и�����-  H�E�H�U�H�M�H�E�H��H��H�	@������H��ЉE��}� u_H��     H�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��и�����  H�EȋU��P,H�EȋPH�Eȋ@ЉE�H�EȋP,H�Eȋ@ �ЋE�ЉE��    I��H��������H���H�E�H�E��    �    H��I��H��s������H��ЋU�H�Eȋ@ H�M��	��H�M���H��:������H��ЉE��E�    �E�    �   �E���Hc�H�E�H�H�E��E�;�l���}~H�E��@a��ta�E���Hc�H��p���H�H�E���   H��H��I��H�%s������H��ЋE���Hc�H��p���H�H��H�H;������H��ЃE����E��}�?�e�����H�E�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��ЋE�H�Đ   [A_]���UH��AWSH��`��H�����I��      L�H�}�H�u�H�U�H�M�D�E�H�E�H�E�H�Eغ�   �    H��I��H��s������H���H�E�H��H��;������H���H��H�E�H��H��I��H�.v������H����E�    �"H�U؋E�H����uH�U؋E�H�� �E��}�_~�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉEп    I��H��������H���H�E�H�EȺ    �    H��I��H��s������H��ЋU�H�E��@ H�M��	��H�Mȉ�H��:������H��ЉEă}� t!H�E�H��I��H���������H��ЋE���  �E�    �$�E���Hc�H�E�H�H�E�H�E��@a��t�E��}�?~���H�E��@a���G  �}�?�=  �U�H�E؉PsH�E��@a��E���H�E؈PbH�U�H�E�H��H��H��<������H���H�U؉BkH�E؋@k���uOH�E�H��H�\�������H�<I�߸    H�f�������H���H�E�H��I��H���������H��и   ��   �E���@��t$H�E؋@kH�U�H�M�H�Ή�H��>������H���H�M�H�E຀   H��H��I��H�%s������H��ЋU�H�E��@ H�M��	��H�Mȉ�H��:������H��ЉEĐH�E�H��I��H���������H��и    �JH�E�H��I��H���������H���H�E�H��H���������H�<I�߸    H�f�������H��Ҹ����H��`[A_]���UH��AWSH��P��H�����I���      Lۉ}�H�u�H�U��    I��H��������H���H�E��E�    �E��E��E������E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E��E܋E�;E���   �}� tV�E�H�U����H�U�H��H�¾   H��:������H��ЉẼ}� t#H�E�H��I��H���������H��и�����?  �E�H�U����H�U�H��H�¾   H��:������H��ЉẼ}� t#H�E�H��I��H���������H��и������   �E��E�E��E��E�   H�E��@�����E�    ��U�E�EȋE�H��    H�E�HЋ �E�E�H��    H�E�H��     �}��uL�E�H�U����H�U�H��H�¾   H��:������H��ЉE̐H�E�H��I��H���������H��ЋE��6�E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��Y���H��P[A_]���UH��AWSH��   ��H�����I�d�      L�H��h����   I��H��������H���H�E�H�E�H�E�H�E�H   H�E�H��h���H�E�H��H��I��H��n������H���H�U�H�E�H��H��I��H��q������H��п   I��H��������H���H�E�H�E��   �    H��I��H��s������H���H��p���H�E�H�E��   �    H��I��H��s������H���H�E��@   H�E��     H�U�H�E�H��H��H��?������H��ЉE�}� t<H�E�H��I��H���������H���H�E�H��I��H���������H��и    ��  H�E�H�U�H�M�H�E�H��H��H�	@������H��ЉE��}� u<H�E�H��I��H���������H���H�E�H��I��H���������H��и�����d  H�E��U��P,H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE��    I��H��������H���H�E�H�E��    �    H��I��H��s������H��ЋU�H�E��@ H�M��	��H�M���H��:������H��ЉE�}� tSH�E�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��ЋE��l  �E�    �   �E������E���Hc�H�E�H�H�E�H�E��@a��t!H�E�H�U�H��H��H�<������H��ЉE�}� u9H�E��@a �U�H�E��@ H�M��	��H�M���H��:������H��ЉE�}� ��E��}�?�k����}� tPH�E�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��ЋE��uH�E��@kH�U�H�M�H�Ή�H�B\������H��ЉE�H�E�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��ЋE�H�Đ   [A_]���UH��H����H�5����I��      Lމ}�E�E��}� u�E��   �E����rH��     H�H��     H�����UH��H����H�����I���      L�H�}��   H�E�H���r�����UH��AWH����H�����I�i�      L�H��     H�H�U�H��     H�    H��       �    H�M�   �    H��I��H��s������H��ѐH��A_]���UH��AWSH��P��H�����I��      Lۉ}��u��}� u
�    ��  H��     H�H=�   v%H���������H�<I�߸    H�f�������H��ҐH��       ���u�H��       ��PH��       ��E����E�E�%�  ��t�E��E�    �E�    �E�    �}� t�E��   �E�   �K  �}��  �=  H��     H�H�E�H�E�    �E�    �  H�E؋@����   H�E؋@9E���   H�E�H�H�E؋@��H�H�E�H�E؋@+E���H�E؉PH�E؋P�E��H�E؉PH�E�H�E�H��     H�H�E��E�    �mH�E؋@��tH�E��E��WH�E�H�E�H�E�H�E�H�E�H�@H�PH�E�H�PH�E��@   H�E�H�U�H�H�E��U��PH�E�H�U�H�P�E���!�}��   ~��H�E��E��}��   ������E�   ���}� ��   H��     H�H�E��E�    �~H�E؋@��tH�E��E��hH�E�H�E��E��H��b������H���H�E�H�E�H�U�H��E��E���H�E��PH�E��U��P�E���+E���H�E��PH�E�H�@   ��}��   �u���H��       �    H��     H�H�PH��     H�H�E�H��P[A_]���UH��SH��(��H�����I���      L�H�}�H�}� ��  �H��       ���u�H��       ��PH��       �H�E�H�E�H��     H�H�E��E�    �M  H�E�H� H9E�tH�E��E��2  H�E�H�E�H��     H�H�P�H��     H�H�E؋@��uH�E�H��H�Pc������H����   H�E؋@��uH�E�H�@H�E�H�E�H�@H�P�H�E�H�PH�E�H�@H��tH�E؋@����   H�E�H�@H��uRH�E�H� H��H�Pc������H���H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    ��}��   �������H��       �    ��H��([]���UH��AWH��H��L�����I���      M�H�}��u�H�E�    �E�    H�}� u�E��   ��H�d������I� ���8  �H��       A� ��u�H��       A� �PH��       A� H��     I� H�E�H�E�H�E��E�    �   H�E�H� H9E�t
H�E��   H�E�H�E��E�   H�E��P�E��=   v@H��     I� �U�H�E�H��H��������I�< M�Ǹ    I�f�������M�A����H�E�H� H�E�H�E��P�E��H�E��P�E��}��   �X���H��       A�     �}� u�E��   ��H�d������I� ���H�E�H��HA_]���UH��H�� ��H�����I��      L�H�}�H�u��E�    H�E�H�E��   H�E�� ��H�E��@9�sH�E��P#H�E��@9�rH�E��@#    H�E�f�   H�E�H�PH�E��@#��H�H�E�H�PH�E�H�PH�U�H�U�H�R� �H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  �E��}��E����E�����UH��H�� ��H�����I��      L�H�}�H�u��E�    H�E�H�E�H�E��@'�PH�E��P'H�E��P'H�E��@9�rH�E��@'   �H�E��P#H�E��@'9�r�H�E��@'�P�H�E��P'�JH�E�H�PH�E��@'��H�H�E�H�PH�E�H�PH�E�H�HH�M���H�E��@'�PH�E��P'�E��}�~��E�����UH��AWSH��0��H�����I�3�      L�H�}�H���������H�H� H�E�H�E�H�E�H�E�H��I��H�
y������H��ЉE�H�E�H��I��H�
y������H��ЉE؋U܋E��=   ~
������   H�E�� </uH�E��E�H�HE�H�m�H�E�� </tH�E�H�E�H�PH�U�� /�H�E�H�U�H�E�H��H��I��H�.v������H���H�E�H��I��H�
y������H��Љ�HE�H�m�H�E�� </u	H�E��  �H�E�H�E��  �    H��0[A_]���UH��AWSH����H�����I��      L�H���������H�H� H��I��H�
y������H��Ѓ�w
�    �   H���������H�H� H�E�H�E�H��I��H�
y������H��Љ�HE��H�E�H�P�H�U��  H�E�� </u�H���������H�H� H��I��H�
y������H��Ѓ�vH�E��  �    H��[A_]���UH��AWSH��0��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
�    ��  H�E�H��I��H�
y������H��ЉE�E�H�H�P�H�E�H�� </u�E�H�H�P�H�E�H��  �}� 
�    �  �}���   H�E�H��� <:u%H�U�H�E�H��H��I��H�.v������H����K  H�<�������H�<I��H���������H���H��H�E�H��H��I��H�.v������H���H�E�H��I��H�
y������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H�.v������H����   H�<�������H�<I��H���������H���H��H�E�H��H��I��H�.v������H���H�E�H��I��H�
y������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H�.v������H���H�E�H��0[A_]���UH��H����H�����I���      L�H�}�H�E�H�E�H�}� u�    �+�E�    �H�E�� </u�E�H�E�H�E�� ��u�E�����UH��AWSH��0��H�����I�J�      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
������   H�E�H��I��H�
y������H��ЉE�E�H�HE�H�m��H�E�� </tH�m�H�E�� ��t�E�P��U�����H�E�H�U�H�E�H��H��I��H�.v������H���H�E��  �    H��0[A_]���UH��H��8��H�����I�e�      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �CH�E�H�PH�U�� ���E�H�E�H�PH�U�� ���E�E�+E�E�}� u�}� t
�m��}� u��E�����UH��H��8��H�����I�ό      L�H�}�H�uЉŰẺE�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M����E��P��U���u�H�E�����UH��H�� ��H�����I�X�      L�H�}���U��E�E��E�H�E�H�E��H�E�H�PH�U��U��m��}� u�H�E�����UH��AWSH��0��H�����I��      L�H�}�H�u�H�E�H�E�H�E�H�E��E�    H�E�H�PH�U�� ����I��H�>�������H��ЉE�H�E�H�PH�U�� ����I��H�>�������H��ЉEԋE�+EԉE܃}� u�}� t뗋E�H��0[A_]���UH��AWSH����H�����I�8�      L�H�}�H�u�H�E�H��I��H�
y������H��Љ�H�E�H�H�E�H��H��I��H�.v������H���H�E�H��[A_]���UH��H�� ��H�����I���      L�H�}�u�H�E�H�E��H�E�� ��9E�uH�E��H�E�H�E�� ��u۸    ����UH��H�� ��H�����I�`�      L�H�}�H�u�H�E�H�E�H�E�H�E��3H�E��H�E�� 8�u!H�E�� ��H�E�� ��Ѕ�u�    �'H�E�H�PH�U��H�E�H�PH�U�� 8�t����������UH��H��0��H�����I�Ɖ      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E��  H�E�����UH��AWH��(��H�����I�I�      L�H�}؉uԋU��҉Uԃ}� uOH�U�H��I��H�
y������H��҉�H�E�H���   H�E�� ��tH�E�� ��9E�u	H�E��   H�E�H�E؃�H��űE�i��E�H�E�H�E��H�E�H�E� ������H�E� ��!�%������u%H�E� 3E䍐����H�E� 3E���!�%������t�H�E�H�E��H�E�H�E�� ��tH�E�� ��9E�u�H�E�H��(A_]���UH��H��@��H�����I� �      L�H�}�H�u�H�U�H�U�H�U������   H�U�H�������   H�E�    H�E�    H�E�    H�E�    �H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�t�H�E�H+E��'H�U����H�Uȉ�H��H��v������H���H+E�����UH��H����H�����I��      L�H�}�H�E�H�E��H�E�H�E�� ��u�H�E�H+E�����UH��AWSH��@��H�����I���      L�H�}�H�u��U�H�E�H�E�H�E�H�E��E�    �kH�E�H�PH�U�� ����I��H�>�������H��ЉE�H�E�H�PH�U�� ����I��H�>�������H��ЉEԋE�+EԉE܃}� u�}� t
�m��}� u��E�H��@[A_]���UH��H��(��H�����I�օ      L�H�}�H�u��U�H�E�H�E�H�E�H�E��}� u)������2H�E�H�PH�U��H�E�H�PH�U�� 8�u�m��}� u����E�����UH��H��8��H�����I�V�      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �!H�U�H�BH�E�H�E�H�HH�M����E��E�9E�w�H�E��  �E�����UH��AWH����H�����I�ׄ      L�H�}�H�u�H�M�H�U�H��H��I��H��w������H��҉�HE�H�E�� ��tH�E���    H��A_]���UH��AWH��(��H�����I�e�      L�H�}؉u�H�U�H��I��H�
y������H��҉E��U�H�E�H�H�E��E�    �H�E�� ��9E�uH�E��H�m��E��E�9E�wڸ    H��(A_]���UH��H��0��H�����I�ԃ      L�H�}�H�u�H�E�H� H�E�H�}� u�    �vH�E�H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u,�}� u
H�E�    �H�E�H���  H�E�H�U�H�H�E���}� u������UH��H��@��H�����I��      L�H�}�H�u�H�E�H�E�H�E�    H�E�    H�E�    H�E�    H�E�� ��u
�    ��   H�E�H��� ��u+�H�E�H�E��H�E�� 8�t�H�E�H+E��   H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�u�H�E�H+E�����UH��H��8��H�����I��      L�H�}�H�u�H�U�H�}� uH�E�H� H�E�H�}� u
�    ��   �H�E�H�PH�U�� ���E�H�E�H�E��
�E�;E�u��H�E�H�PH�U�� ���E��}� uۃ}� uH�E�H�     �    �   H�E�H��H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u4�}� u
H�E�    �H�E�H��H�E�H�E��  H�E�H�U�H�H�E���}� u������UH��H����H�����I���      L�H�}�H�u�H�u�H�M�H��       H�H��H�~������H�������UH��AWSH�� ��H�����I�S�      L�H�}�H�u�H�E�H��I��H�
y������H��ЉE��2�U�H�M�H�E�H��H��I��H��r������H��Ѕ�uH�E��H�E�H�E�� ��uø    H�� [A_]���UH��AWSH�� ��H�����I��      L�H�}�H�E�H��I��H�
y������H��Ѓ��E�E��I��H��������H���H�E�H�}� u�    �$�U�H�M�H�E�H��H��I��H�%s������H��АH�� [A_]���UH��H��8��H�����I�      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��U�H�E�H�H�E�H�E�H;E�v[H�E�H;E�sQH�E�H�E��E�HE��H�m�H�m�H�E��H�E��H�E�H;E�u��'H�U�H�BH�E�H�E�H�HH�M���H�E�H;E�u�H�E�����UH��AWH����H�����I�Z~      L�H�}�H�u�H�M�H�U�H��H��I��H��u������H���H��A_]���UH��AWH����H�����I�~      Lډ}�H�@�������H�<I�׸    H�f�������H�������UH��H����H�����I��}      L؉}��U���H���������H�Hc��������t�E� �E�����UH��H����H�����I�a}      L؉}��U���H���������H�Hc��������t�m� �E�����UH��AWSH��0��H�����I�	}      L�H�}ȉuĉU��M��U�H�E�H��H�P�������H�<I�߸    I�f�������I�A��H�E�H��I��H���������H���H�E�H�E� �E�H�E� 9E�u��H��0[A_]���UH��AWSH�� ��H�����I�g|      L�H�}�H�u�H�E�� ��u�    �LH�E�� <wuH�E�H��I��H���������H���H�U�H�E�H��H��I��H��1������H���H�E�H�E�H�� [A_]���UH��AWH����H�����I��{      L�H�}�H�U�H��I��H�D3������H���H��A_]���UH��AWH����H�����I��{      L�H�}�H�U�H��I��H�]2������H���H��A_]���UH��AWH����H�����I�<{      L؉}�H�u�H�M��U�H�Ή�I��H��3������H���H��A_]���UH��AWSH�� ��H�����I��z      L�H�}�H�}� u������VH�E�H��I��H��5������H��ЉE�H�E؋@��u+H���������H�H��E�H�։�I��H��3������H��ЋE�H�� [A_]���UH��AWH����H�����I�Qz      L؉}�H�u�H�M��U�H�Ή�I��H���������H���H��A_]���UH��AWH����H�����I��y      L�H�}�H�U�H��I��H�	�������H���H��A_]���UH��AWSH��@��H�����I��y      L�H�}ȉu�H�U�H�}� u	H�E��  H�E�H�E�H�E�H�E��E�    H�E�H��I��H��5������H��ЉEԃ}����   H�E��@��u7�}�u�}� ~+H���������H�H��E�H�։�I��H��3������H��Ѓ}�
tk�E�;E�}E�}�u�}� ~H�E�H;E�vH�m��m��:�}��^���H�E�H�PH�U�UԈ�E��D����}�u�}� ~�m���E��)�������}�~	H�E��  ��Eԉ�H�E�H�E�H��@[A_]���UH��AWSH�� ��H�����I�Wx      L�H�}�H�u�H�}� u�    �^�E�    �2�E�Hc�H�E�H�� ��H�U�H�։�I��H���������H��ЃE�H�E�H��I��H�
y������H��ЋU�9�w��E�H�� [A_]���UH��AWH��(��H�����I��w      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I��7������I�A��H��(A_]���UH��AWH��(��H�����I�Ww      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I�b8������I�A��H��(A_]���UH��AWH����H�����I��v      L�H�}�H�U�H��I��H��^������H���H��A_]���UH��AWH����H�����I��v      L�H�}�H�U�H��I��H�5:������H��ҐH��A_]���UH��AWH��(��H�����I�cv      L�H�}�H�u��U܋U�H�u�H�M�H��I��H�9������H���H��(A_]���UH��H����H�����I�v      L�H�}�H�}� u������!H�E��P#H�E���+  9�r�������    ����UH��AWH����H�����I��u      L�H�}�H�U�H��I��H��9������H���H��A_]���UH��AWSH��`  ��H�����I�bu      L�H������H������H�������E�    �E�    �  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H��������H���	E�}���  �E�H��    H��i  H�H��i  H�>��H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E��E�H������H�։�I��H���������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�}� t(H������H�E�H��H��I��H���������H����O  H������H��H�h�������H�<I��H���������H����   H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E�H�������E�H�։�I��H�_�������H���H������H������H��H��I��H���������H����w  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������
   H��H��I��H���������H���H������H������H��H��I��H���������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������   H��H��I��H���������H���H������H������H��H��I��H���������H����  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�EȾ   H��fHn�I��H���������H���H������H������H��H��I��H���������H����]  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eк
   H��H��I��H�1�������H���H������H������H��H��I��H���������H����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ
   H��H��I��H���������H���H������H������H��H��I��H���������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ   H��H��I��H���������H���H������H������H��H��I��H���������H����G  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�E�   H��fHn�I��H���������H���H������H������H��H��I��H���������H����   H������H�ƿ%   I��H���������H��ЋE�Hc�H������H�� ��H������H�։�I��H���������H����4�E�Hc�H������H�� ��H������H�։�I��H���������H��ЃE��E�Hc�H������H�� ��������    H��`  [A_]���UH��H����H�����I��l      L؉��E��E�    �E��S��%wa��H��    H��b  H�H��b  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I�(l      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��H�� ��H�����I�Bk      L�H�}�H�u�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E�����UH��AWSH��  ��H�����I��j      L�H������H������H��x����E�    H������H�E�f�E�  �E� �E�    �/  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H��������H���	E܃}���  �E�H��    H�Na  H�H�Ca  H�>��H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E��E�H�U�H�E�H��H��H���������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H�}� t'H�U�H�E�H��H��H���������H���H�E��e  H�E�H�`�������H�4H��H���������H���H�E��7  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E�H�������E�H�։�I��H�_�������H���H������H�E�H��H��H���������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������
   H��H��I��H���������H���H������H�E�H��H��H���������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������   H��H��I��H���������H���H������H�E�H��H��H���������H���H�E��3  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�E��   H��fHn�I��H���������H���H������H�E�H��H��H���������H���H�E��x  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�E��
   H��H��I��H�1�������H���H������H�E�H��H��H���������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ
   H��H��I��H���������H���H������H�E�H��H��H���������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ   H��H��I��H���������H���H������H�E�H��H��H���������H���H�E��e  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�Eо   H��fHn�I��H���������H���H������H�E�H��H��H���������H���H�E��   H�E�H�g�������H�4H��H���������H���H�E�fǅ����  �E�Hc�H������H�� ������H������H�E�H��H��H���������H���H�E��8�E�Hc�H������H�� �E�H�U�H�E�H��H��H���������H���H�E��E��E�Hc�H������H�� �������H�E��  H�U�H������H)�H��H�Ā  [A_]���UH��H����H�����I�b      L؉��E��E�    �E��S��%wa��H��    H��Y  H�H��Y  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I�Ra      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H��������L��Љ�<�����<���Hc�H�����H��  ��<���H���   A_]���UH��AWH���   ��L�����I�Q`      M�H����������H�����H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H����������H�����H��M��H���������L��Љ�<�����<���H���   A_]���UH��AWSH��0��H�����I�f_      L�H�}؉u�H�U�H�M��}�   v
�    �   H�U�H�E�H��H��       H�<I��H��������H��ЉE�}���  ~�   �I�E�E�}� ~:�U�H�E�H��       H�4H��I��H�%s������H��ЋE�Hc�H�E�H��  �E�H��0[A_]���UH��AWH����H�����I��^      L؉}�H���������H�H�
�U�H�Ή�I��H���������H���H��A_]���UH��AWSH�� ��H�����I�1^      L�H�}�H�}� tj�E�    �?H���������H�H��E�Hc�H�E�H�� ��H�։�I��H���������H��ЃE�H�E�H��I��H�
y������H��ЋU�9�w���H�� [A_]���UH��AWH���   ��L�����I��]      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I��\      M�H��8���H��0���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�H�`�������I�<M�׸    H�f�������L�������UH��AWH����H�����I��[      L�H�}�H�U�H��I��H���������H��ҐH��A_]���UH��AWH��(��H�����I��[      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H�?�������H��Ѹ    H��(A_]���UH��AWH��(��H�����I�E[      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H�?�������H����H�E�H�E�� < tH�E�H   H9E�sH�E�� <
u�H�E��  H�E�H;E�����H��(A_]���UH��AWSH��0��H�����I��Z      L�H�}�H�uЉỦM�H��      H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H�?�������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H��      H�H�E�H��      �0H��      �D �}�u-�U�H�E�    H��I��H��������H���H�U�H��   �}�u+�U�H�E�    H��I��H�2�������H��Љ�H�EЉ�[�}�u,�U�H�E�    H��I��H�2�������H��Љ�H�E�f��)�U�H�E�    H��I��H�2�������H��Љ�H�EЈ�    H��0[A_]���UH��AWSH��0��H�����I��X      L�H�}�H�uЉỦM�H��     H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H�?�������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H��     H�H�E�H��     �0H��     �D �}�u'H�E�H��I��H��������H����Z�H�E�� �+�}�u%H�E�H��I��H��������H���fH~�H�U�H��    H��0[A_]���UH��SH��8��H�����I��W      L�H�}�H�u�H�U��E�    �E�    ��  �E�    �E�Hc�H�E�H�� ������%��  �E��E�Hc�H�E�H�� ������lu�E��E�   �E�Hc�H�E�H�� ����H���������H���	E�}��o  �E�H��    H�pP  H�H�eP  H�>��H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H�H�������H�����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H���������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�O�������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�O�������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��������H����?  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�O�������H�����   H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�O�������H����jH�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��������H������E��E�Hc�H�E�H�� ��������E�H��8[]���UH��H����H�����I�hS      L؉��E��E�    �E��S��%wa��H��    H�_M  H�H�TM  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��R      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H�0�������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I��Q      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H�0�������L��Љ�<�����<���H���   A_]���UH��H����H�����I��P      L؉}�H�u�H�}� u������w�}��u������jH�E��@#��tH�E��@#�P�H�E��P#H�E��@#H�U��J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U���E�����UH��AWSH����H�����I�)P      L�H���������H�H� H��I��H��5������H��ЉE�}��t+H���������H�H��E�H�։�I��H��3������H��ЋE�H��[A_]���UH��AWH��(��H�����I��O      L�H�}�H�u�H�U�H�h�������H�<I�ϸ    H�f�������H�������UH��H����H�����I�FO      L�H�}��	   H�E�H���r�����UH��SH����H�����I�O      L�H�}�H�}� u.H��     H�<H���������H���H��     H��H�E�H��H���������H���H�E�H��[]���UH��AWSH��0��H�����I��N      L�H�}�H�u�H�E�H�z�������H�4H��I��H���������H���H�E�H�}� u
������   �E�    H�E�H��I��H�
y������H��ЉE܃}�`~	�E�   �$H�E�H�P+H�E�H��H��I��H�.v������H���H�E��@���H�E��PH�E�H��I��H� �������H��ЋE�H��0[A_]���UH��H��0��H�����I��M      L؉}�H�u�H�E�H�E��E܉E��E�    �}� y,H�E�H�PH�U�� -�}�   �u�E�����E���E��؉E�H�E�H�E�M�Hc�Hi�gfffH�� ��������)�����)��ʉЍH0H�E�H�PH�U�ʈ�E�Hc�Hi�gfffH�� ����)ЉE�}� u��}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWSH��@��H�����I�KL      L�H�}�H�u��U�H�}� u#H�E�H�E�H�E�H�PH�U�� 0H�E��  �  H�E�H�E؋E�Hc�H�E�H�H�E��3H�E؃��E�H�m��}�	~�7   ��0   �U��H�m���H�E�H�E�H;E�wËE�Hc�H�E�H��  H�E�H�E��E�    �8H�E�� <0uH�E��"H�U�H�E�H��H��I��H�.v������H�����E��E�;E�|�H�E�H�E�H�E�H��I��H�
y������H��Љ�H�E؋E�H�U�)Љ�H�M�H�E�HȾ    H��I��H��s������H���H��@[A_]���UH��AWH����H�����I��J      L؉}�U�    ��I��H�d������H���H��A_]���UH��AWH����H�����I��J      L؉}�u�U��U��I��H��������H���H��A_]���UH��AWH����H�����I�;J      L�H�}�H�U�H��I��H�7g������H��ҐH��A_]���UH��AWH����H�����I��I      L�H�}�u�M�H�U��H��I��H�8i������H���H��A_]���UH��H����H�����I��I      L؉}�u�E��}�E��E��}�ЉE��}� x�E���y�E����E��E�+E�E��!�}� y�E���~�E����E��U��E�ЉE�H�E�����UH��H�� ��H�����I�I      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H�� ��H�����I�lH      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H��H��H�����I��G      L�H�}�H�u��U�H�E�H�E�H�E�H�PH�U�� ���E�E���H���������H�H������ ��uǃ}�-u�E�   H�E�H�PH�U�� ���E��"�E�    �}�+uH�E�H�PH�U�� ���E�}� t�}�u9�}�0u3H�E�� <xtH�E�� <XuH�E�H��� ���E�H�E��E�   �}� u�}�0u�   ��
   �E��}� t	H��   ������H�E�E�Hc�H�E�H�H��H�ЉE؋E�Hc�H�E�H�H��H�E�}� t�}� ~�E�)E�H�E��]�H�E�    �E�    �E���H���������H�H��������t�m�0�[�E���H���������H�H���������5  �E���H���������H�H��������t�7   ��W   )E�E�;E���   �}� ��   �}� tgH�E�H;E�|H�E�H;E�u0�E�;E�~(�E�����H�E�   �H���������H�� �����   �E�   �E�H�H�U�H��H�E��E�H�H)E��eH�E�H;E�H�E�H;E�u-�E�;E�~%�E�����H�E����H���������H�� �����$�E�   �E�H�H�U�H��H�E��E�H�HE���H�E�H�PH�U�� ���E��y������H�}� t�}� t
H�E�H���H�E�H�U�H�H�E�����UH��AWH����H�����I��D      L�H�}�H�M�
   �    H��I��H�2�������H���H��A_]���UH��AWH����H�����I�9D      L�H�}�H�M�
   �    H��I��H�2�������H���H��A_]���UH��AWAVAUATSH����H�����I��C      L�H�}�H�uȉU�L�eп    L��L�`� �؉���H���������H�H������ ��uЃ�-u�   L��L�`� �����+uL��L�`� �؃}� t�}�u-��0u(A�$<xt	A�$<XuI�D$� ��I���E�   �}� u��0u�   ��
   �EċE�Hc������    H��I�ǋE�Hc������    H��H�Љ�A�    A�    ����H���������H�H��������t��0�T����H���������H�H��������tz����H���������H�H��������t�7   ��W   )�;]�}GE��x
M9�wM9�u��9�~A������A�   �E�H�L��Hc�I�L��L�`� ���;������E��yA�����H���������H�� "   �	����tI��H�}� tE��tI�D$��H�E�H�U�H�L��H��[A\A]A^A_]���UH��H����H�����I��A      L؉}��   �   ���r����UH��AWSH����H�����I�`A      L�H�}�H�E�H�}�������H�4H��I��H��u������H��Ѕ�uH���������H�H� ��    H��[A_]���UH��AUATSH�� ��H�����I��@      L�H�}�H�u�H�8     ��E�L�e�H�]�E�,$L��L�`��H��H�XD�(�m��}� uې�H�� [A\A]]���UH��H��8��H�����I�q@      L�H�}�H�u�H�U�H�8     ��E�H�E�H�E�H�E�H�E�H�E�H�E�H�E�� ���E�H�E�H�PH�U�H�U���H�E�H�PH�U�H�U���H�E�H�PH�U��U���m��}� u�������UH��SH��H��H�����I��?      L�H�}�H�u�H�8     ��E�H�E�H+E��EȋE�9E���  �E�����EȺ    ��E��EȋU�H�E�H�H�E�H�E�H�E�H�E�H�E�E�H�H��H��H�E�H�H�E�H�E�H;E�sjH�0     H�H�U�H�E�H��H���щEă}� u/�E�H�H��HE�H�U�H�E�H��H��H��������H�����  �}� y�E�H�HE���  �H�E�H;E���   H�0     H�H�U�H�E�H��H���щEă}� u)�E�H�HE�H�U�H�E�H��H��H��������H���뢃}� ��   H�E�H;E�uA�E�H�HE�H�U�H�M�H�E�H��H��H���������H��ЋE�H�HE�H�E�H�E��M���H�U�H�E�H��H��H��������H��ЋE�H�H��HE��E�H�HE���   �E�H�H��HE�����H�E�H;E���   H�E�H+E�H��H�E�H+E�H9�|4�E�Hc�H�E�H�H�E�H��H��H�1�������H���H�E�H�E������H�U�H�E�H��H��H�1�������H��ЋE�Hc�H�E�H�H�E������E�H�H��HE�H�U�H�M�H�E�H��H��H���������H��ЋE�H�H��HE�H�E�H�E������H��H[]���UH��H�� ��H�����I��<      L�H�}��u�U�H�M�H�0     H�U�H��U�H�8     ��U��U���H�U�H�H�U�H��H��H�1�������H��А����UH��AWH����H�����I�N<      L�H�}�H���������H�<I�׸    H�f�������H��Ѹ����H��A_]���UH��H��@��H�����I��;      L�H�}�H�u�H�U�H�U��H�E�H�U����H���������H�Hc���҃� ��u��E�    H�U���҃�+t��-u�E�   H�E�H�����������E��E�    �E�    �E�    �;�M�H�����������Y�H�U���҃�0�*��X��E�H�E��E�H�U����H���������H�Hc���҃���u�H�U����.uuH�E��?�M�H�����������Y�H�U���҃�0�*��X��E�H�E��E��E�H�U����H���������H�Hc���҃���u��U�)U�}� uH���������f���  �}� t�E�H���������f(fW��E�H�U����etH�U����E��   �E�    H�E�H�U���҃�+t��-u�E�   H�E��E�    �%�M܉����҉�H�U���҃�0ʉU�H�E�H�U����H���������H�Hc���҃���u��}� t�U�)U���U�U�}����|	�}�   ~H�����������   H�����������E��E�E܃}� yF�]��A�E܃���t&�}� y�E��^E��E���E��YE��E��}��E��Y��E��}� u�H�}� tH�E�H�U�H��E�����UH��H����H�����I��8      L؉}�H�E�   �E�    �H�U�H��H��H�H�H�E��E��E�;E�|�H�E�����UH��AWSH��@��H�����I�]8      L��E�H�}��u�H�}� u	H�E��  H�E�H�E�H���������f��f/E�v,H�E�H�PH�U�� -�E�H���������f(fW��E��E�H���������f/s�E��H,�H�E��/�E�H�����������\��H,�H�E�H�       �H1E�H�E�H�E�H�E�H��x�H*��H��H���H	��H*��X��M��\�f(��EȋE���H�5�������H���H��x�H*��H��H���H	��H*��X��YE�H���������f/s�H,�H�E��*H�����������\��H,�H�E�H�       �H1E�H�E�H�E�H�M�H�U�H�E�H���������H�43H��I�߸    I���������I�A��H�E�H��@[A_]���UH��AWH����H�����I�s6      L�H�}�H�U�    H��I��H� �������H���H��A_]���UH��AWH����H�����I�#6      L�H�}�H�u�H�M�H�U�H��H��I��H� �������H����Z�H��A_]���UH��AWH��(��H�����I��5      L�H�}�H�u�H�M�H�U�H��H��I��H� �������H����E��E�H��(A_]���UH��H����H�����I�m5      L؉}��E����3E�)�����UH��H��@��H�����I�95      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�    H�}� y>H�E�H�PH�U�� -H�       �H9E�uH��������H�E�H�E��H�E�H��H�E�H�E�H�E�H�M�H�gfffffffH��H��H��H��H��?H)�H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U��ʈH�M�H�gfffffffH��H��H��H��H��?H)�H��H�E�H�}� u�H�}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U߈H�E�H;E�w�H�E�����UH��AWH��8��H�����I��3      L�H�}�H�uЉU�H�U�H�U�H�}� yH�U�H�JH�M��-H�]�H�U�H�U��}�u$H�M�H�u�   H��I��H���������H����H�M�H�U�H��H��H���������H���H�E�H��8A_]���UH��H��0��H�����I�3      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E�H�M�H���������H��H��H��H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U�ʈH�E�H���������H��H��H��H�E�H�}� u�H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWH��8��H�����I�2      L�H�}�H�uЉU�H�U�H�U�H�U�H�U��}�u$H�u�H�M�   H��I��H���������H����H�M�H�U�H��H��H���������H���H�E�H��8A_]���UH��H����H�����I��1      L؉}������UH����H�����I�`1      Lظ   ]���UH��H����H�����I�51      L�H�}��    ����UH��H����H�����I�1      L�H�}�H���������H�H� ����UH��H����H�����I��0      L�H�}�H���������H�H� ����UH��H�� ��H�����I��0      L�H�}��u�H�U�H�M�    ����UH����H�����I�Z0      Lظ    ]���UH��H����H�����I�/0      L��E�H���������f������UH��H����H�����I��/      L��E�H���������f������UH��H����H�����I��/      L��E��}�H���������f������UH��H����H�����I��/      L��E�H�}�H���������f������UH��H����H�����I�D/      L��E��M�H���������f������UH��H��(��H�����I�/      L��E��M��E��U��U��E��E��E������������������������������]��E�����UH��H����H�����I��.      L��E����E����]��E�����UH��H����H�����I�].      L��E�H���������f������UH��H����H�����I�$.      L��E�H���������f������UH��H����H�����I��-      L��E�H� �������f������UH��H����H�����I��-      L��E�H����������E��E�����UH��H����H�����I�n-      L��E�H��������f������UH��H����H�����I�5-      L��E�H��������f������UH��H����H�����I��,      L��E�H� �������f������UH��H����H�����I��,      L��E�H�(�������f������UH��AWH����H�����I��,      L��E��E�H�0�������H�f(�fHn�I��H���������H���H��A_]���UH��H����H�����I�),      L؉}�H�u�    ����UH��AWH����H�����I��+      Lډ}�H�u�H�8�������H�<I�׸    H�f�������H�������UH��AWH��(��H�����I��+      Lى}�H�u�H�U�H�I�������H�<I�ϸ    H�f�������H�������UH��AWSH�� ��H�����I�H+      L�H�}�H�]�������H�<I�߸    H�f�������H����E�    �.�E�H�H��    H�E�HЋ ��I��H�d�������H��ЃE��}�?~̸����H�� [A_]���UH��AWH����H�����I��*      L�H�}�u�H�n�������H�<I�׸    H�f�������H�����f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f�                                                                    ~ � � � � � � � � ~             ~ � � � � � � � � ~                 l � � � � | 8                   8 | � | 8                   < < � � �   <                < ~ � � ~   <                      < <              � � � � � � � � � � � � � � � �           < f B B f <           � � � � � � � � � � � � � � � �        2 x � � � � x             < f f f f <  ~               ? 3 ? 0 0 0 0 p � �              c  c c c c g � � �               � < � < �             � � � � � � � � � � �               > � >                  < ~    ~ <                f f f f f f f   f f              � � � {                | � ` 8 l � � l 8  � |                       � � � �              < ~    ~ <  ~              < ~                           ~ <                      �                         0 ` � ` 0                         � � � �                       ( l � l (                      8 8 | | � �                   � � | | 8 8                                                 < < <                  f f f $                             l l � l l l � l l           | � � � |   � � |               � �   0 ` � �             8 l l 8 v � � � � v           0 0 0 `                             0 0 0 0 0 0               0         0                   f < � < f                         ~                                    0                     �                                                           0 ` � �             8 l � � � � � � l 8              8 x       ~             | �    0 ` � � �             | �   <    � |               < l � �                 � � � � �    � |             8 ` � � � � � � � |             � �     0 0 0 0             | � � � | � � � � |             | � � � ~     x                                                       0                  0 ` 0                      ~     ~                     ` 0      0 `             | � �                       | � � � � � � � |              8 l � � � � � � �             � f f f | f f f f �             < f � � � � � � f <             � l f f f f f f l �             � f b h x h ` b f �             � f b h x h ` ` ` �             < f � � � � � � f :             � � � � � � � � � �             <         <                   � � � x             � f f l x x l f f �             � ` ` ` ` ` ` b f �             � � � � � � � � � �             � � � � � � � � � �             | � � � � � � � � |             � f f f | ` ` ` ` �             | � � � � � � � � |           � f f f | l f f f �             | � � ` 8   � � |             ~ ~ Z       <             � � � � � � � � � |             � � � � � � � l 8              � � � � � � � � � l             � � l | 8 8 | l � �             f f f f <     <             � � �   0 ` � � �             < 0 0 0 0 0 0 0 0 <               � � � p 8                 <         <          8 l �                                                   �       0                                     x  | � � � v             � ` ` x l f f f f |                   | � � � � � |                < l � � � � v                   | � � � � � |              6 2 0 x 0 0 0 0 x                   v � � � � � |  � x       � ` ` l v f f f f �                 8      <                        f f <       � ` ` f l x x l f �             8         <                   � � � � � � �                   � f f f f f f                   | � � � � � |                   � f f f f f | ` ` �             v � � � � � |                � v f ` ` ` �                   | � ` 8  � |              0 0 � 0 0 0 0 6                    � � � � � � v                   � � � � � l 8                   � � � � � � l                   � l 8 8 8 l �                   � � � � � � ~   �             � �  0 ` � �                 p                                        p         p                       v �                        8 l � � � �                               ��� ��� ~~~                                 uuu ��� ��� ���                                 ��� ��� ��� ��� ;;;                          ��� ��� ~~~ ��� ���                         ��� ��� ���     ��� ���                         ��� ���      ��� ��� ppp                 @@@ ��� ���         III ��� ���                 ��� ��� ��� ��� ��� ��� ��� ���                 ��� ���                 zzz ��� ���         ``` ��� ���                     ��� ���         ��� ��� MMM                     ��� ��� bbb     ��� ���                         ||| ��� ���      ��Cw Simples editor File  Open  Save  Close  Exit  Help    Y���������������Y�������Y�������Z�������Z�������Z�������Z�������Z�������Z�������Z�������Z�������Z�������Z�������Z�������Y�������BitMAP error
 Not suport BitMAP 4-bit Not suport BitMAP > 8-bit ____ none
 File name    KIB MiB GiB ./ File %s %lf            �@      �A      0AEntrada maior que o limite
 Erro ao criar o arquivo "%s"
       Error ao criar o arquivo "%s", atingio o limite de arquivos na entrada de directorio
   Panic: __malloc, sem espaco na tabela de alocacao
      panic: realoc sem espaco, %lx size = %d %d
 PWD strerrorr
      (((((�AAAAAABBBBBB                                �Dubug: %s %x %x
        (null)  ����������������������]����������������������d�������d������������������������������������������������������������������������������������ �������Қ��������������6�������6�������T���������������������������������������o���������������������������������������������������������������������������������������K�������]�����������������������x���������������]�������������������������������������������������������������������������������T���������������f�����������������������o�������(null) %        ��������Þ������N�������	���������������_�������������������������������������������������������������������������������������������������������������Ȣ������y�������*�������ۤ������ۤ������*�������`�������`�������`�������`�������E�������`�������`�������`�������`�������`�������`�������`�������`�������`�������`�������!�������3�������`�������W�������N�������`�������3�������`�������`�������`�������`�������`�������`�������`�������`�������`�������*�������`�������<�������`�������`�������E�������panic: sscanf()
        ����������������������k�������װ�������������C�������C��������������������������������������������������������������������������������������������������������������������������������������������������������������ֲ������������������������������������������������������������������������������������Ĳ��������������������߲�������������Ĳ������������������������������������������������������������������������������������Ͳ��������������������ֲ������panic: freopen()
 r+ PWD call system funtion error. 
                 $@       �        %lu.%lu                �              �C                                                                        �_�
�@panic: signal()
 panic: sigaction()
 panic: setjmp()  panic: longjmp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �C �     �     �    U �   �C �   8U �   �C �      �   �C �      �   �C �   �4 �   �C �   D �                                   x3 �   |3 �   �3 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  zR x�  ,      @����   E�CG����B�A�       $   L   �����    E�CG����B�A�   t   �����   E�CG��  ,   �   U���   E�CG���B�A�          �   <����    E�C�� $   �   ����   E�CE��A�   $     �����    E�CG����B�A�$   4  &����    E�CG����B�A�(   \  �����   E�CG����B�A�   (   �  C���j   E�CG��W�B�A�       �  �����    E�CE���� (   �  ���   E�CG���B�A�         ����    E�CE���� (   (  �����   E�CG��q�B�A�   $   T  ����   E�CG����B�A�   |  ����9    E�Cp�     �  ����+    E�Cb�     �  �����    E�C��     �  l����   E�CE����      ���I    E�C@�        7���u    E�CE�f�A�(   D  �����   E�CG����B�A�   (   p  >����   E�CG����B�A�   $   �  �����    E�CG����B�A�,   �  ����2   E�CG���B�A�       (   �  ����D   E�CG��1�B�A�   $      �����    E�CG����B�A�(   H  :����   E�CG����B�A�   ,   t  ����   E�CG����B�A�       ,   �  ����   E�CG���B�A�       (   �  �����   E�CG��s�B�A�   $      �����    E�CG����B�A�(   (  ����   E�CG��
�B�A�   $   T  �����    E�CG����B�A�$   |  #���   E�CF��A�   (   �  ����   E�CG����B�A�   $   �  �����    E�CG����B�A�(   �  >���5   E�CG��"�B�A�   $   $  G���k    E�CG��X�B�A�   L  �����    E�C��    l  .����    E�C��    �  ����X    E�CO� ,   �  
���l   E�CG��Y�B�A�       ,   �  F���6   E�CG��#�B�A�       (     L���D   E�CG��1�B�A�   (   8  d ��q   E�CG��^�B�A�   (   d  ����   E�CG����B�A�   (   �  m���   E�CG����B�A�   (   �  ���Z   E�CG��G�B�A�      �  ��   E�C�      	���    E�C��    (  �	���    E�C��     H  
��p    E�CF�`�A�$   l  ]
���    E�CG����B�A�$   �  ��r    E�CG��_�B�A�(   �  f��   E�CG��	�B�A�   $   �  V���   E�CF���A�       	  ����    E�CE���A�    4	  ����    E�CE���A�   X	  *���    E�C��    x	  ���A    E�Cx�      �	  	��i    E�C`�        �	  N��U    E�CL�    �	  ���U    E�CL�    �	  ���i    E�C`�    
  ��g    E�C^�    <
  H���    E�C�� $   \
  ���   E�CE�{�A�      �
  q��9    E�Cp�  $   �
  ����    E�CG����B�A�   �
  K��^    E�CU� (   �
  ���   E�CG���B�A�   (     r���   E�CG����B�A�   (   D  ��]   E�CG��J�B�A�   (   p  A��   E�CG��l�B�A�   (   �  ���D   E�CJ��.�B�A�   (   �  �%��:   E�CG��'�B�A�   $   �  �&��    E�CG����B�A�     �'���    E�C��    <  F(���    E�C�� (   \  �(���   E�CJ����B�A�   (   �  �,��i   E�CG��V�B�A�   (   �  �/��H   E�CG��5�B�A�   (   �  2��e   E�CJ��O�B�A�        O6��a    E�CX�    ,  �6��9    E�Cp�      L  �6���    E�CF�w�A�(   p  7��'   E�CG���B�A�   $   �  :��   E�CE���A�   $   �  �;���   E�CF���A�      �  Z=��    E�C��      :>���    E�C�� (   ,  �>��O   E�CG��<�B�A�   $   X  !@���    E�CG����B�A�(   �  �@��C   E�CG��0�B�A�      �  �B��k    E�Cb� $   �  GC���    E�CG����B�A�   �  D���    E�C��      }D��w    E�Cn�    4  �D��b    E�CY� $   T  E���    E�CG����B�A�$   |  �E��z    E�CG��g�B�A�   �  �E��a    E�CX�    �  <F���    E�C��    �  �F��{    E�Cr� $     G��+   E�CF��A�      ,  H��6   E�C-�   L  *I��L    E�CC� $   l  VI���    E�CG����B�A�   �  �I���    E�Cw�    �  VJ��}    E�Ct� $   �  �J��r    E�CF�b�A�    $   �  �J���    E�CF���A�       $  hK���    E�C��    D  L��3   E�C*�   d  M��7   E�C.�   �  /N��W    E�CN� $   �  fN���    E�CG����B�A�$   �  �N���    E�CG����B�A�   �  NO���    E�C�� $     �O��V    E�CF�F�A�       <  P��P    E�CF�       \  NP��U    E�CL�    |  �P��U    E�CL� $   �  �P���    E�CG����B�A�$   �  2Q���    E�CG����B�A�$   �  �Q��K    E�CF�{�A�     $     �Q��K    E�CF�{�A�     $   <  �Q��S    E�CF�C�A�    $   d  R���    E�CG����B�A�$   �  �R��S    E�CF�C�A�    $   �  �R��K    E�CF�{�A�     ,   �  �R��[   E�CG��H�B�A�       $     �S���    E�CG����B�A�$   4  vT��]    E�CF�M�A�    $   \  �T��]    E�CF�M�A�    $   �  �T��K    E�CF�{�A�     $   �  U��L    E�CF�|�A�     $   �  'U��Y    E�CF�I�A�       �  XU��Y    E�CP� $     �U��K    E�CF�{�A�     (   D  �U���   E�CJ��{�B�A�       p  ^���    E�C��     $   �  �^���    E�CI���A�       �  b_��l    E�Cc� (   �  �_���   E�CJ����B�A�         Wh���    E�C��     $   ,  �h��   E�CI���A�    $   T  �i���    E�CI���A�    $   |  {j���    E�CG����B�A�$   �  ,k��\    E�CF�L�A�    $   �  `k���    E�CG����B�A�$   �  �k���    E�CI���A�         �l���    E�CI�    $   <  ,m��L    E�CF�|�A�         d  Pm��e    E�CF�U�A�    �  �m���    E�CF���A�(   �  n���   E�CG����B�A�   (   �  �o��=   E�CG��*�B�A�   $     �p��\   E�CE�M�A�      ,  �t���    E�C�� $   L  Vu���    E�CI���A�    $   t  v���    E�CI���A�       �  �v���    E�C�� $   �  xw���    E�CG��z�B�A�   �  �w��Y    E�CF�         x��9    E�Cp�  $   $  /x���    E�CE�q�A�    $   L  �x���    E�CG����B�A�   t  Wy��G   E�C>�,   �  ~z��u   E�CG��b�B�A�       $   �  �{��M    E�CF�}�A�     $   �  �{��O    E�CF��A�     $     |��L    E�CF�|�A�     $   <  3|��S    E�CF�C�A�       d  ^|���    E�C�    �  �|���    E�C��    �  P}���    E�C��    �  �}��2   E�C)�$   �  ���U    E�CF�E�A�    $     ���U    E�CF�E�A�    4   4  F���L   E�CM�����-�B�B�B�B�A�      l  Z���7    E�C       $   �  q���w    E�CG��d�B�A�(   �  ����{    E�CI���d�B�B�A�   �  ����    E�C�� $      �����   E�CE���A�       (  g����    E�Cx�     $   L  ć��\    E�CF�L�A�       t  ����5   E�C,�   �  ���_    E�CV� ,   �  L����   E�CG����B�A�       $   �  ���P    E�CF�@�A�    $     /���Z    E�CF�J�A�    $   4  a���^    E�CF�N�A�       \  ����4    E�Ck�     |  ����v   E�Cm�$   �  ����    E�CF���A�       �  �����    E�C�� $   �  a����    E�CF���A�         ΐ��*    E�Ca�     ,  ؐ��'    E�C^�     L  ߐ��/    E�Cf�     l  ���;    E�Cr�     �  	���;    E�Cr�     �  $���:    E�Cq�     �  >���'    E�C^�     �  E���9    E�Cp�       ^���9    E�Cp�     ,  w���<    E�Cs�     L  ����=    E�Ct�     l  ����>    E�Cu�     �  Α��n    E�Ce�    �  ���;    E�Cr�     �  7���9    E�Cp�     �  P���9    E�Cp�        i���9    E�Cp�     ,   ����D    E�C{�     L   ����9    E�Cp�     l   ����9    E�Cp�     �   ؒ��9    E�Cp�     �   ���9    E�Cp�  $   �   
���a    E�CF�Q�A�       �   C���2    E�Ci�     !  U���T    E�CF�   0!  ����X    E�CF�$   L!  ɓ���    E�CG����B�A�   t!  <���T    E�CF�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    GCC: (Ubuntu 9.3.0-17ubuntu1~20.04) 9.3.0                                        �                    �                  @ �                 p@ �                 �@ �                 �@ �                  ` �                                     ��                     ��_ cole _             ��                )        �           ^         �           0    ��                7    ��                @     <"  �   �       G      h2 �           L      j2 �           Q      y2 �           V      2 �           [      �2 �           `      �2 �           e      �2 �           j      �2 �           o    ��                u    ��                �    ��                �    ��                G       3 �           L      .3 �           Q      F3 �           �    ��                �    ��                �    ��                �     EI  �         �    ��                �    ��                G      `3 �           �    ��                �     �@ �          �    �@ �          �     �@ �          G      e3 �           �    ��                �    ��                G      k3 �           �    ��                �    ��                     �@ �           
     A �               �@ �          �     i  �   �      !    l  �   �      V      �3 �           [      �3 �           `      �3 �           e      �3 �           j      �3 �           &     �3 �           +     �3 �           0     �3 �           6   ��                =   ��                G      �3 �           L      �3 �           Q      �3 �           �   ��                C     A �          G      H4 �           L      �4 �           S   ��                Z   ��                G      �4 �           a   ��                j   ��                s   ��                |   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                   ��                   ��                    (A �          $   ��                -   ��                6   ��                @   ��                J   ��                G      �4 �           U   ��                ]   ��                g   ��                q   ��                G      �5 �           y   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �    ��  �   �       G      �5 �           �   ��                �   ��                �    c�  �   �       G      �7 �           L      �7 �           �   ��                   ��                   ��                    @A �             ��                �   ��                �   ��                #   ��                G      �9 �           ,   ��                5   ��                ?    ��  �   e       v    �  �   �       T    ��  �   �      I    @A �          S    c�  �   =      Z    @B �          �    ��  �   �       6   ��                7   ��                d   ��                m   ��                w   ��                G      �; �           �   ��                �    @C �   `       �   ��                G      �; �           �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                G      �; �              ��                    �C �              �C �              x�  �   {           ��  �   �       &    �  �   �      *   ��                G      �; �           3   ��                G      < �           L      < �           Q       < �           <   ��                C    � �   _       G      8< �           L      @< �           Q      P< �           V      0< �           N   ��                U   ��                ^   ��                h   ��                n   ��                u   ��                |   ��                }   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                G      X< �           �   ��                �   ��                �   ��                G      `< �           �   ��                G      h< �           �   ��                G      p< �           �   ��                G      x< �           �   ��                G      �< �           �   ��                G      �< �           �   ��                G      �< �           �   ��                G      �< �           �   ��                G      �< �           �   ��                �   ��                G      �< �           L      �< �              ��                G      �< �           L      �< �                ��                    p@ �           #    � �   T       +    y�  �         �    ��  �   \       >    �O  �         H    9-  �   �       S    ��  �   {       Z    n �   9       ^    � �   ;       c     �   �       j    2  �   �       z    �?  �   �       ~    ��  �   7      _    ��  �   �       �    �C �          �    ��  �   �      �    ��  �   �       �      �               �(  �   �       �      �           �    ^�  �   P       �    P �   �       �     U �          �    F�  �   �       �    �  �   �       �    �C �          �    ��  �   �      �    )�  �   U       �    [9  �   u       �    �  �   w       �    � �   9       �    8U �          �    h �   9           �
 �   ^           `2 �              �%  �             � �   �       P    ��  �   �       "    ��  �   [      (    x�  �   :      4    ��  �   �       D    �g  �   q      �
    y�  �   �       P    ��  �   w       W    �5  �   �           fM  �   �      f    �<  �   �      n    l�  �   L       u    + �   v      �    0�  �   �       |    ��  �   U       �     �   \       �    X�  �   Y       �    ��  �   M       �    h�  �   K       +
    �C �          �     M �          �    �]  �   �       �    L6  �   �      �    � �   <       �    ��  �   �       �    �F  �   �      �    ~�  �   L      �    ��  �   G      �    �C �          �    �o  �         �    X�  �   ]          ^)  �   �       K    �L �   4           ��  �   K       $       �           )    %*  �   �      2    �9  �   �      9     ` �           B    �n  �   Z      L    }�  �   �       R    dz  �   A       Y    ƹ  �   �       e    q@  �   2      l    &b  �   6      s    �x  �   �       {    ��  �   2      �    �C �          �    ��  �   �       �    �r  �   �       �    ��  �   �       �    �E  �   �       �    I �   �       �    ��  �   O       �    p �   5      �    HK  �         J	     D �   �       �    �z  �   i       �    �^  �   l      �    �	 �   P       ^    7�  �   �       �    :[  �   5      �    �y  �   �       �    )�  �   z       �    ��  �   �      o     � �               X�  �   �           ��  �   Y           �T  �         +    ��  �   9       :    Z�  �   �      C     �   �      <    / �   9       H    �C �          N       �          ~
    �@ �           W    (U �          ]       �           d    �C �          m     � �           s    �  �   �       z    �~  �   9       �    !|  �   g       �
    � �   D       �	     �   '       �      �   >       �    m �   T       �    �  �   V       �    ��  �   �       �    c{  �   U       �    �'  �         �    ^ �   n       �    �  �   }       �    '  �   �       �    n�  �   �       �    5 �   9       �     M �          �    s�  �   S       	    �+  �   j      	    ��  �   k       	    ��  �         
    �@ �           '	    ��  �   W       .	    ��  �   H      9	    ��  �   �       �    �D �          @	    ��  �   �       G	    �  �   �       S	    ��  �          ^	    J�  �          i	    � �   X       s	    x  �   �       z	    ��  �   �       �    �C  �   D      �	    ��  �   ]       �	    �4 �          �	    4�  �   D      �	    0U �          �	    o}  �   �      �	    ��  �   �       �	    �D �          �	    ��  �   �       "
       �           �	    �  �   9       �	    � �   ;       �	    �  �   b       �	    �C �          �	    "#  �   �      �	    ��  �   K       �	    � �   *       �	    �S  �   �       	
    ��  �   K       
    8�  �   �           / �   /       
    �s  �   r        
       �           '
    �C �          �    W�  �   �       �    � �   a       2
    ��  �         �
    &�  �   S       ;
    �5  �   +       �    Bv  �   �      I
    �q  �   �       Q
    "�  �   l       E    &t  �         [
    �  �   �       �
    � �   9       b
    9  �   I       h
    b^  �   X       q
    ��  �   e      }
    �@ �           �
     �   9       �
    d�  �   K       �    �  �         �
    �-  �         �
    ?
 �   Z       �
    D�  �   6      �
    y �   9       �
    � �   �       �
    ; �   2       Q    ��  �   �       �
    �C �          �
    I�  �   i      �
    ��  �   �       �
    q  �   �       �
    ��  �   '      '    N�  �   �       !
       �           �     D �          �
    �  �   S       �
    ]r  �   p       �
     0 �   @      �
    N   �               i�  �   C          � �   :            �  �   u      &    ��  �   �       ,    �  �   ]       3    �U  �   �      ?    D �          n     � �           H    o\  �   k       O    ��  �   \      W    ��  �   L       ^    ��  �   Y       f    �\  �   �       �       �           p    J�  �   �       z    ��  �   7           D �          �    ZZ  �   �       �    _�  �   a       �    ��  �   U       -    T4  �         �    ��  �   �       �    �D �          A    �/  �   �      �    �{  �   i       �    ^ �   ;       �    M�  �   3      �    `   �   �      �    /  �   �       �    z�  �   L       �       �           �    �  �   U       �    [5  �   9       �    �|  �   �           �N  �   �            �   '       �       �               �  �   ^       (    ��  �   �       *    �
 �   4       .    ��  �   a       5    
�  �   �       ;    @ �   9       @    �  �   +      J    \e  �   D      W    � �   =       ]    ��  �   �      f    ��  �   r       n    {  �   U       z    '�  �   L           .�  �   O       lib/setup.asm HEADER_MAGIC HEADER_FLAGS header crt0.c editor.c gravar .LC0 .LC1 .LC2 .LC3 .LC4 .LC5 .LC6 .LC7 gui.c font8x16.c window.c bmp.c font.c border.c editbox.c editbox_refresh mouse.c menubox.c obj.c objm foc message.c dialog.c button.c listbox.c file_data file_type file_unidade attr .LC8 .LC9 .LC10 file.c cfs.c alloc_spin_lock pipe.c path.c memcmp.c memcpy.c memset.c strcasecmp.c strcat.c strchr.c strcmp.c strcpy.c strcspn.c string.c strlen.c strncasecmp.c strncmp.c strncpy.c strpbrk.c strrchr.c strsep.c strspn.c strtok.c last.1481 strstr.c strdup.c memmove.c strcoll.c strerror.c ctype.c tolower.c toupper.c stdio.c fopen.c fclose.c fflush.c fputc.c fgetc.c fgets.c fputs.c fread.c fwrite.c remove.c rewind.c fseek.c feof.c ftell.c vfprintf.c vf vsprintf.c vsnprintf.c sn_buf putchar.c sscanf.c perror.c vfscanf.c character _buf.1638 fvalue _buf.1650 ungetc.c getchar.c freopen.c tmpnam.c _tmpnam rename.c itoa.c i2hex.c malloc.c calloc.c free.c realloc.c lldiv.c strtol.c atoi.c atol.c strtoul.c exit.c getenv.c qsort.c qscmp qses qsexc qstexc qs1 system.c strtod.c ftoa.c _precision atof.c strtof.c strtold.c abs.c ltoa.c utoa.c srand.c errno.c gmtime.c localtime.c strftime.c clock.c math.c pow.c sqrt.c atan.c acos.c asin.c floor.c ceil.c exp.c locale.c signal.c setjmp.c _GLOBAL_OFFSET_TABLE_ longjmp read_directory_blk menumotor drawstring strcpy log sqrt setjmp clean_blk_enter put strtok_r stdout vsprintf ungetc pwd_ptr argv strerror utoa_r __m_i memmove __tm __realloc_r atol __window_puts getenv ceil errno floor strtold _infinity loop qsort fgets file_update file_read_block m_file_list memcpy __window_clear BitMAP2 perror ltoa_r tolower system feof malloc remove fs_directory msg_read __window_putchar ldexp vsnprintf m_edit strtoul itoa __pipe__ stdgetc_r update_directory_entry _drawline fflush argc drawrect BitMAP eh_frame stdputc_r upath tell_r strncasecmp border button write_r strtol user rename flush_r strrchr update_editbox utoa calloc strtod fmouse rewind_r dialogbox atof update_objs seek_r strcat read_directory_entry debug_o fseek obj_focprocess __free_block_r open_dir ftoa stdin font8x16 __m_c _start obj_list __end strstr write_blk get_file_name atan2 signal strcoll strncmp write_sector draw_char_transparent pow strncpy put_pixel strcasecmp log10 _BLK_ realloc drawchar path_count open_file_r strtok remove_blk memcmp sscanf getfilename file_close pipe_write sigaction read_r file_write_block fread _ctype open_file addr search_blk_null strdup save fopen sysgettmpnam localtime memset pwd main ftell srand init_process fclose getchar close_r __data ptr_mouse2 __free_r update_window getkeyw _vsputs_r strcmp color msg_init remove_file __bss atan fgetc drawchar_trans strtof strcspn asin ltoa setlocale stderr create_file strsep getkey __malloc_r fputc open_r A__ call_function getpathname strftime i2hex lldiv fwrite obj_process __window getmsg vfscanf rewind freopen msg_write pipe_read exit pipe_r register_obj __block_r atoi __heap_r ptr_obj assert_fn gmtime strspn ctr0 drawstring_trans strlen __code toupper wcl filename_cmp submenubox clock read_super_block abs strchr fputs acos strchrnul file_listbox frexp vfprintf strpbrk read_sector free setpath  .symtab .strtab .shstrtab .text .data .got .got.plt .data.rel.local .bss .eh_frame .comment                                                                                     �                                       !                �                                          '              @ �    @     p                              ,             p@ �   p@                                  5             �@ �   �@                                   E             �@ �   �@     @                             J              ` �    P      0                             T      0                �     *                                                   0�     h.      
   �                 	                      ��     �                                                   �     ]                                                                                                                                                                                                                                                                                                                                                                                                                              BM��     6  (   �  �            �  �                                                          	         
  
     
      


  

              
 
                            $ (	 $ , # , ( 6 % ' 1 +# 9& -$ *$ 7) 85 $ " &$ *! """ &&& *** ... +(% 7,% ;3* 444 <<< ;88 ./1 # G F( H7 O3 G9) G<6 S9( g; YF pM YF+ WI9 MG6 mT4 we3 ~b CCC MMM KGG VMG [TK UUU \\\ ]YV PPQ hYH h]U oXK ldY xjX xjN ddd lkk utu }}} xxy yqh \_f ?@6 �q2 �f# �v[ �rR �zj �}u �{i �qP ��9 ��8 ̗< ��T ��Y ��S ��V ��k ��x ��s ��h ��z ��p ��h ��s ɜV ʧY ժQ �W Ǜf ɛv ɨi ϭp �` ��t ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ʳ� ƻ� 붃 �Ʋ �׾ ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �� nde                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 Q -
  .J                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     QQiJ .                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            M N� p                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
����j-                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ������J.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ������M.                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����߿                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �����lP                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         $B\ CJ  J+                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 SO B��M
 -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ]B:��+  
  *                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            3]��Y  *K                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               B:1��VVM 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             XX��Yw2    
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            6o��Ww[6KK+  
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �n�yT66T-*  +
                                                                                                                                                                                                                                                                                                                                                                                                                                                             'I<a748b�z g                                                                                                                                                                                                                                                                                                                                                                                                                                                                    I'R=:b��7BN%                                                                                                                                                                                                                                                                                                                                                                                                                                                                          O:3V��7B +'                                                                                                                                                                                                                                                                                                                                                                                                                                                                          OO3��3\ N                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     834��4@8*I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    978��18Y37EE                                                                                                                                                                                                                                                                                                                                                                                                                                                                      b:V��2y13<$MD                                                                                                                                                                                                                                                                                                                                                                                                                                                                      cZ��ZW8V\e                                                                                                                                                                                                                                                                                                                                                              ���r  "                                                                                                  J <<=1��V:Z                                                                                                                                                                                                                                                                                                                                                            .�����k                                                                                                  	*<<=��ZV11:                                                                                                                                                                                                                                                                                                                                                            �����                                                                                                     9X\1���                                                                                                                                                                                                                                                                                                                                                             �����p    $                                                                                                  a4Bn��3a \                                                                                                                                                                                                                                                                                                                                                            R����� R3  $                                                                                                  BB:Y�{< <P                                                                                                                                                                                                                                                                                                                                                             ���J\9"                                                                                                  B\V��W B]N0                                                                                                                                                                                                                                                                                                                                                            ...MK- ��\ 9$                                                                                                ]b1��6WL,S)K*                                                                                                                                                                                                                                                                                                                                                            i   r�z779                                                                                                \b��V[TNNM EE'                                                                                                                                                                                                                                                                                                                                                                
��Y:@:9                                                                                  e)B922Y2��<O+                                                                                                                                                                                                                                                                                                                                                                                  

T��c81B                                                                                  %e=226��V<+                                                                                                                                                                                                                                                                                                                                                                                 

4c�cc=                                                                                  		 E466��c$-                                                                                                                                                                                                                                                                                                                                                                                  
::��c:7                                                                                  		) <a2��`:X                                                                                                                                                                                                                                                                                                                                                                                
1YY��X                                                                                 3Xc1��c2aB+                                                                                                                                                                                                                                                                                                                                                                               84cY�zB                                                                                OBVy�4:BB")                                                                                                                                                                                                                                                                                                                                                                               a3��:8                                                                                		Z1Z2W�Tc4=0)                                                                                                                                                                                                                                                                                                                                                                            
   nX\��X                                                                                		Zc2Y��TWcYN                                                                                                                                                                                                                                                                                                                                                                                    O9X�\:\B                                                                                %.N$2Yy��4Z8                                                                                                                                                                                                                                                                                                                                                                                    R��X89B"                                                                                ')jV2 2::V                                                                                                                                                                                                                                                                                                                                                                                    M9:��1a4 "                                                                                EnY��Z\:\                                                                                                                                                                                                                                                                                                                                                                                    <\b�y@87<                                                                                ,A9:8��48cB                                                                                                                                                                                                                                                                                                                                                                                    %%*, X:��ab$                                                                                  \9Y:6��X=\ M                                                                                                                                                                                                                                                                                                                                                                                     DI =8:Y��@O                                                                                 =]1T��c6\< *                                                                                                                                                                                                                                                                                                                                                                                    II\11cc�cX9                                                                                MM\T{�v]= =-                                                                                                                                                                                                                                                                                                                                                                                     EFE 48y`z�b9                                                                                k$8��wWz]33                                                                                                                                                                                                                                                                                                                                                                                         91��T`['                                                                )M$Vc2]��(g%%%%                                                                                                                                                                                                                                                                                                                                                                                      X1n�{[['                                                                I	9cTX�n](;%%%%                                                                                                                                                                                                                                                                                                                                                                                      9X��W[                                                                E08V66WĎX                                                                                                                                                                                                                                                                                                                                                                                      71Xc��T,"'                                                                '08VTT��Y:9                                                                                                                                                                                                                                                                                                                                                                                      <38YY�w9                                                                 !(5^66Y��3@7$                                                                                                                                                                                                                                                                                                                                                                                       B22��b9                                                                 ;(=X2w��TZ3@Z9                                                                                                                                                                                                                                                                                                                                                                                    		    b9\2��Y1@"                                                                =>4=1]��cY79$AN                                                                                                                                                                                                                                                                                                                                                                                    		    ]O 3Xy�{48,                                                                \===4��Vy@ 9jS                                                                                                                                                                                                                                                                                                                                                                                            ��YT@:<                                                        *   KK+C\b��n9,E	&F&&	                                                                                                                                                                                                                                                                                                                                                                                    T��c:8<                                                        J    pM B�o$��7M%F&&%''))%		                                                                                                                                                                                                                                                                                                                                                                                           6w�cn49                                                         J p- �����l?iGG('                                                                                                                                                                                                                                                                                                                                                                                             TT��cX                                                         
  .  �������RN,G''***                                                                                                                                                                                                                                                                                                                                                                             6`Y��\                                                        *   .��������<n:1166W[111113!!                                                                                                                                                                                                                                                                                                                                                                                        6Tc`�zB                                                        +
 jP���������B:11T6W`::8488                                                                                                                                                                                                                                                                                                                                                                                        `2:4��B=                                                        k   ���������8`��}~xx~[WWWWWTTT6621111                                                                                                                                                                                                                                                                                                                                                                                w61V\��\                                                        r QP���������4w²����������{wYWTT::==                                                                                                                                                                                                                                                                                                                                                                                    0\4c�`W[X3%                      -L9$ X4�� �������3=W������������������������~|xxv[T6666TWUU248:983  )::::88771111((((!!!!%%%%%%%%%%%%		                                                                                                                                                                                                                                                                    < ::��WT:X&                      .-/0" 794=��a������B:�}���������������������������������{ycXX:89B]a
)+)3333787$77$4211;;((!!!%%%%%%%%%%%		                                                                                                                                                                                                                                                                    ::T��6c4'                             //]7=X8=��a\9$qǕ +)GG<O::WWW[TW`dw��������������������������������~~~}v[[```UUUUUUUUUU222222&&%%%%&&%&&&&&&&  ''%%&&&&111      !!!!!!!!######55                                                                                                                                                                                                                                                                    *"1Y6`�{V:$E                          .PM ,+9=3o�naBX<) 	RE91:WVT6[[WWT:TT[[[[[`vv~~�������������������������������{{wwc^UU666>>2''&&DDFFDDD&&&&&%%&&DDDD11111433333377!!!!!!!!######55                                                                                                                                                                                                                                                                    F%+<8TV��1cb$                      9BB��on="] #ItI%D&%%HO;$< 777379:UUUUUUU^W[xx{�������������������������������~}x``[[[[[[WWUWW[[v77778888		      ####1155                                                                                                                                                                                                                                                                    'E,92ZY��VO                      EP+*C79��zB<-RM)%fD&&%!! 89UUUUUUUUUUWWWUWWuu[[uv|~|���������������������������������|xv[WUZVV@@@884444;;>>           ####1155                                                                                                                                                                                                                                                                    EF]3cc�cZ:                          M/7B��]\3=<EIE?.I%%DFFFFFF&   DDDDDDDDDD'5;;>>511]]X6226Xww���������������������������������~~|xvuuu[[[[????$?$?DDDD!!!!%%%%%%&&&&DDDDDD&&%%                                                                                                                                                                                                                                                                    e&e:ybz�b:                          gSR�Ǖ���3\9m<)t#-%&kefFHF&DF))))IIJ+fFDDDDDDfII)))HOOO=>5166662222```[T666`vxx|����������������������������������dd__CC$$$$((FFFF!!!!%%%%%%&&&&DDDDDD&&%%                                                                                                                                                                                                                                                                    B@��48:  *                ) 
J""����ɑ\  3<77798:::VVVVW[``{���������������������������������~|||xTT6TWWWT6622:T:2221155+)I) ** ,  +                                                                                                                                                                                                                                                            73o�y18
 	                 + O<m������b95<    778844446:TWWWWWUUUUvv|~����������������������������������`[T:TWYY2212>=<<)+)e-JM  
*                                                                                                                                                                                                                                                            B��2:33	                 S\=]z�����$<!!!!;;;;;;;;


	################&&%%%%%%&DFFFFEE\XO==8877:V_`w����������������������������������~||vv[6W61!g&&pqpR 
                                                                                                                                                                                                                                                            BY��:83                 =4nX������,""!!!!;;;;;;;;


	################DDD&&&%%%%548::@@@77777U[uu[[uv~~������������������������������w`11O(&����r                                                                                                                                                                                                                                                               /3 XY�{T214                AT:n��\�ŉA   /(((((((((((;;;;;;DDDDDDDD'DDDDD((,00,DD&% 
+HHFF(("599CCCC__W[x{��������������������U22>>������P+                                                                                                                                                                                                                                                              B:4��Y21:                 Ry12��cX\r  	(((((((((((;;;;;;DDDDDDDD&&&''D''				%%))----++FD((HHOO$$UUWWUUW[uuuuu|�����������U62n������  
                                                                                                                                                                                                                                                            P$a:Ð[2T                 C\b1z��6W1X 9EF'*	  %%!!((((''''''''''((''2221111111111111<<+"?$$Z@@9871((((EFFD%<<<9 HHhH>><<maa$m�����+P                                                                                                                                                                                                                                                              geXc��{6:                 $O B��y6�T128�bn))*	'  %%!!((((''''''''''((''2211111111111222NOOL<+$+??????99A<<;;55"@@@@8843==H>H;;(FDDD%%00<<9973hhhH>;;=o $B?#����MRk

                                                                                                                                                                                                                                                                        
��V1 9B7%%  #	 %&GS= Z@9W6w��YO'!S6��v &&%%                                                                                                                                                                                                                                                                                                                                                                                                                                                 

X��Y X%%    %%0!9 _@6��w6T5"F!M6��v &&%%                                                                                                                                                                                                                                                                                                                                                                                                                                                 

6n�cb B%%      		78B@��y14:4<E"G6y�v3&&%%                                                                                                                                                                                                                                                                                                                                                                                                                                                 
::��c@7%%  		

"\ ��YVY:OI"0:Y�x3&&%%                                                                                                                                                                                                                                                                                                                                                                                                                                               
1]Y��3\	7�Ĉ99BMP,:V�31%&%%                                                                                                                                                                                                                                                                                                                                                                                                                                               16ncB	yÙ9B8"BB3eT6��31%&%%                                                                                                                                                                                                                                                                                                                                                                                                                                               ]X:��9 !!!! 9@_��y98m)<j<$ e*V8��44%%%                                                                                                                                                                                                                                                                                                                                                                                                                                            
   ]1ac��@!!(! 9CZ��o@=95Re i *V8�44%%%                                                                                                                                                                                                                                                                                                                                                                                                                                                    5] \�n!]]O=@c��dZ <;!) -1{�:T F'                                                                                                                                                                                                                                                                                                                                                                                                                                                    > ��gG("7\=o��_@9 (! *x�cT ''                                                                                                                                                                                                                                                                                                                                                                                                                                                    !99$��"@98B��n C%%''W��: 3')                                                                                                                                                                                                                                                                                                                                                                                                                                                    0\a�OO" <78zÑ 8 %%'' 6��69)                                                                                                                                                                                                                                                                                                                                                                                                                                                    F'-+$!9n ��:]B<"!
	'''"1��68*                                                                                                                                                                                                                                                                                                                                                                                                                                                    %I*AOS 9���Zb8N"  
F'E"4��T33'                                                                                                                                                                                                                                                                                                                                                                                                                                                    DF t#$NM�����b7@@OG&%		E%&I=a�[:                                                                                                                                                                                                                                                                                                                                                                                                                                                    eDP �������c@$ O0&&''	 E'%PX:�`B                                                                                                                                                                                                                                                                                                                                                                                                                                                    b�������                              
�WV 		                                                                                                                                                                                                                                                                                                                                                                                                                                                    p������                              
��VV 		                                                                                                                                                                                                                                                                                                                                                                                                                                                    l�������                              
��VV                                                                                                                                                                                                                                                                                                                                                                                                                                                     ������                              
��WV                                                                                                                                                                                                                                                                                                                                                                                                                                                     �����r                              
�`V                                                                                                                                                                                                                                                                                                                                                                                                                                                      a�                              
{�yV9 *                                                                                                                                                                                                                                                                                                                                                                                                                                                    O<�]9                               
{��VB ,                                                                                                                                                                                                                                                                                                                                                                                                                                                    O$a�\9\                              
{��WX ,                                                                                                                                                                                                                                                                                                                                                                                                                                                     9��9=                                6��:7BL                                                                                                                                                                                                                                                                                                                                                                                                                                                     z�98                                6�V7B/                                                                                                                                                                                                                                                                                                                                                                                                                                                    a�9:1                                4d�c3:,                                                                                                                                                                                                                                                                                                                                                                                                                                                      B�9:                                8W�y7!!                                                                                                                                                                                                                                                                                                                                                                                                                                                      73�X:1                                V:��"                                                                                                                                                                                                                                                                                                                                                                                                                                                      93�n61                                Z4��7"                                                                                                                                                                                                                                                                                                                                                                                                                                                       51��62                                Z4��B"                                                                                                                                                                                                                                                                                                                                                                                                                                                    33z�:4                                Z4��\"                                                                                                                                                                                                                                                                                                                                                                                                                                                    SB]�:8                        7Y�{T2Y                                                                                                                                                                                                                                                                                                                                                                                                                                                    MO\�X8                        7V��T2X                                                                                                                                                                                                                                                                                                                                                                                                                                                    LOB�b8                        76��T4:                                                                                                                                                                                                                                                                                                                                                                                                                                                    ,A7�y8                        74��T66                                                                                                                                                                                                                                                                                                                                                                                                                                                    /< ��8                        3:��T:1                                                                                                                                                                                                                                                                                                                                                                                                                                                    Nz�8                        9Vy�[:1                                                                                                                                                                                                                                                                                                                                                                                                                                                    M< a�:                        \Xc�wV1                                                                                                                                                                                                                                                                                                                                                                                                                                                    SO \�:                        ]XY�Z1                                                                                                                                                                                                                                                                                                                                                                                                                                                    <03 �\                         :1��::                                                                                                                                                                                                                                                                                                                                                                                                                                                    /,73�n!                         :4��V:                                                                                                                                                                                                                                                                                                                                                                                                                                                    +77y�"                        48�V:                                                                                                                                                                                                                                                                                                                                                                                                                                                      0"39X�! 
                        (1=c�_:                                                                                                                                                                                                                                                                                                                                                                                                                                                      / =4�! 
                        G=W�w:                                                                                                                                                                                                                                                                                                                                                                                                                                                    < 9�< 
                        G9V��:                                                                                                                                                                                                                                                                                                                                                                                                                                                    / 33�i<                         P33W��:                                                                                                                                                                                                                                                                                                                                                                                                                                                    033�pO                        e3Y��:                                                                                                                                                                                                                                                                                                                                                                                                                     RN  N - * J
 * ,N -Q M   * P  *
P
l    ��BAQ eJ *   P . P .-  .   
$n��_9G%&*  --  PJ 
,*+ 
  -iQ  J   N  .K   -.  M M  M  kM J+ + p  .J                                                                                                                                                                                                                                                                                                                                                     - .  *Q
  KrR -p*P P
 +  M-
 j  *�cb  RPM   K*PJ   j  j   
$bB��@]!GF%  P 
N
N-  j* +.M   K -M M
p  K 
j+  
--J+MM .  
P Q  +                                                                                                                                                                                                                                                                                                                                               ir R  j. i  N  K.  
  
   PJP,  . Qj MR�c NS
MM- 
-- JJ P J. i-  Sc9\b(%E  
*-K.K N  J  *J+ M  P  Miii R -J  l ,K Q  iP  P..  +  .j  MQj                                                                                                                                                                                                                                                                                                                                             Q����K
*��
  
-*  q������K+��P ��r   ǿP�B�І<-��k R, k߽l -N�  
��s S@_����=9GG&&*  * �����
   -  ��. , K*P����rp  . ��l, -*������k+ R��N-��j+��p +                                                                                                                                                                                                                                                                                                                                             ��Ŋ�݊ ,��-
  *- J�տ���  M �� P*��  *��p�z��O  P��s -j֋M
ܿ+ k��R y��í��\<%%**  *P�ʔ�޽.    KݗPK i  �އ���K  . ��ki p R�ɽ���r*+p��J��ll��MJ+                                                                                                                                                                                                                                                                                                                                            r��i.�J,-��  -* P�-RMKM, +�� 
 ��M 
p��pJ����$<*ME��q . R Q�
  .ȽJ-���r A�ؙ�c��Q!%&  -,.��J �� *R  j��Q   ��Q.��p J ��qM N P��jN+M . .��Pk��.�� N,                                                                                                                                                                                                                                                                                                                                            K޿ ,Q��J  P��Q M.   JR�  -*  Q��K, ��j  
Q�������  I�ׅ  *K p׾P+ k��k ��� ���n��jGF
QJ ��-,��.M M Q��K    ��RP �֕ J Q�ȅl  i  ��    l K�� ��� ��  
                                                                                                                                                                                                                                                                                                                                            ���  j��Nk  �� k. 
 JQ�P* K -Pi��M.��p . �Ȗ����Kq��MQ*l M֗- ipӖkN���� $��yď��oONrM  �� ..��Q*-RݿM .rl-p�jN��rK
P ��qR  P ���pK p*p j��P���� �� i                                                                                                                                                                                                                                                                                                                                            P��M ��    ��r-MKp  QjߗjN-   J��MP��  ,*��QX�� ��s	, k�, ,Mɿ.�޾�eA��c���؈N"N KJ, .P�ս,
 r��Q  .+N*. q��- N-J �Ҍ  , 
J�� Jj  +��*�Ř�Q��k 
                                                                                                                                                                                                                                                                                                                                            k��P  ��  K����ՕM Jq߾p i K.  ��ǽ��  ,*��j9��\$- ��s	, k�, ,MҾK�Ֆ�e<��_�Ġ�ni0e* ++ J���J .
* ���R *.- - ���lP- * �Ҍ  , 
K�ՆKM J��M��qԇ��i                                                                                                                                                                                                                                                                                                                                             l��R  ��  -�҆��ׅ .r�����l+- ������P   +��r ��$J ��s	, k�, ,ֿi�ǋ�i,��Z����b'E   
J���JPp  +����J P  ���Q*R KP �Ҍ  , 
R����� 
J ��r�pMɖ��Q
                                                                                                                                                                                                                                                                                                                                             R��P ��.   ��ii�
 
r�Ȕ��PJ+ *��*���  -j�@��9$ 
��s	, k�, , �ŊӔ��s��Y���a9-  *���M     p��ܾR   r��l J .  �Ҍ  , 
l�֗q�k  �Ӗ�Q����Q                                                                                                                                                                                                                                                                                                                                              RܿP ��Q,
 ��j��-  �߽ N   .R��Ri��J  .ݗc��9 
��s	, k�, ,���p��p"��byāz9M- , Q��-PK KR 
�Ջ��P, J��Q -
  k
+�Ҍ  , 
��+ *-
+  ���� l����i                                                                                                                                                                                                                                                                                                                                              k׾R  ��   ,��JMQ��.*qܖ JP*K . ��J  ��Q  J �Ə��$+ ��s	, k�, ,jӿݽP��r0��cZ���y". 

-��* N .  ��Pq܊ .�ֽk  P    �Ҍ  , 
�� -- K ��ݾkk���i                                                                                                                                                                                                                                                                                                                                             l��Q  ��-  �� QȿMM,pֽ ,   �� J ��j  K
 �����7+* ��s	, k�, ,q���M��q<��yV�cN$Ii  .P��jMQ��iM k�� ��NK ,�օq ��q** JP�Ҍ  , 
M�� *JM M *���j
���i 
                                                                                                                                                                                                                                                                                                                                            Q��R  ��kPJ�� M�ҽp  ���RJ -. l��*p��k  M

���ڙa< 
��s	, k�, ,q���-Mq��0��b���cAq  iP�Ջ�-��  
K�Ȗ,��kp *q߾M ��,M   +�Ҍ  , 
p��M*JQ K 
��ߊ k ���Q 
                                                                                                                                                                                                                                                                                                                                            +��Җ�Ն  - �ӽ���j  Mi��Ž�� Q-*���ܖ -+*PP�����qž��˭�a Nj֊*M J��� *��IiL�۠�ѬY3E'M  + -�Ř�� 
+��iN-�� K-J�׋���N*P�������,RNj�ӿ���� MP��� . 
���.J                                                                                                                                                                                                                                                                                                                                             -J���ҕ-K  �����q + j������,+k����ʽp 
  l���a�]l�������  lӽM  ��q .��PR<z���� @<g  ,i ���ܽJJM *ֿ  M�� 
p M����* j�������    ������ql J���   ���MQ                                                                                                                                                                                                                                                                                                                                             Qi++J--KP        M
Ri- JJ   J.
K 
,-K  a9�l  PiPiS/mm KM  ,Q,R.KJ))jgB_� c( 
 *j  l P  M K--* MR ,J*MMJ P* ijK**   Q Rk  R
M  J* J JK                                                                                                                                                                                                                                                                                                                                              ,  .Q   M-   -P  J KQ  
+M. 
i-  -     Ji.c8B�O]iM   + P KM 
 ..  
II ]c�cbG(   J JM KJ   P   -  - *+-  .  Q* . N M   R   +   Q *+
 *J-.
                                                                                                                                                                                                                                                                                                                                                  Ki-* J  *Q Ji    
   i-     J  .i, -$S�lk	P)-  *  J P  * I!Y�yb<  N Kj   +    J 
  - *
 K      J .Q+  +
  -P    J
    J                                                                                                                                                                                                                                                                                                                                            .J.  -P  .     ,j*
  -J* N     - K    , J*n����sr)E+GS R . J  p
  +)Ia=n��Y .K   
PK
*-K* K   ,  **,  J Q  i N-PJQkQi.* R      K
                                                                                                                                                                                                                                                                                                                                                 K-   .MJJ  k- Q       KK  -P   JQ 
+   ������M  M  M,   
 
IGbo�bk *,RJ 
M..-      
, KR     *  R   -  ,*      iN  *  K*-  M                                                                                                                                                                                                                                                                                                                                            jP

-  RjP l+-  
 PMjP*. 
 kM   *Qi*+   p+������jsKMggi
 .Q  iMMjQ**MPG <����$(Rk     ii

 , M .   Kp  *P* kP  .KipJR  iMKP
.ilN  -. p +,                                                                                                                                                                                                                                                                                                                                              M    


     
*   


  ,
  PMk���׿ MP            
 e0����m$'            .                          ,              NR           
  
     ..*.+***  
   *,, 
     ,        -*   
 -  
   

 
++ ,K
  ,                                                                                                                                                                                                                                            *     *
  J-,--+
            
-
   -����K  K'0    + 0(������+g' -
                           -K.  *     .           ,.
  ,-.*    
  
*+RPK-


          J
         P
KP   -J   -P*
   
-N-
      
  
J-                                                                                                                                                                                                                                                 JPM         
     **
     ., P. j<$+)           -
*'%������,0        
  
                         Q
.PM
             *         
-*     
*JN          -  KP **-*   
               ,MiM 

     *   .     
                                                                                                                                                                                                                                                
* J**KM.
 JKMQl�������qkK
K+
*,*     -a]EP        *M*  +Eq����b        P*MM--                          , .M        MMM  -        ,
.  +   
-N*Mkq��������piN-.PJ        +           .-  *iK   Q�������qpi-    *M    J*                                                                                                                                                                                                                                              -  -R
   p�����������������Կ�rR. -N  O  ME,,,,,,,,R  ..iQAFr�ʛRj,,,,,,,,K JJ   M                        .  ,-,,,,,,,,KQNK
N            *.* -
 P��������������������Ǖk.,MK  
          ,     Qii�����������������ƕrQM   
                                                                                                                                                                                                                                            ,     Kq�������������������������Խ�-J  *,  
$9BB9 +����������������҅QG'QA���������������טJ  
                        �����������������r  *             +-j���������������������������ǅ.J
- 
K          
MR+ *Q����������������������׾R  KPN                                                                                                                                                                                                                                            *  +-�������������������������������֕j ,  -]XB�\b J+������������������]	0&%'EJ#�����������������                            l�����������������p
.
         
  R, r�������������������������������֗+ 
.
,          ,*k�����������������������������r                                                                                                                                                                                                                                                 iM. P�����������������������������������޽i - o]9zˬ�8aB)M������������������RA		E%'jKt����������������iJN                        l������������������-  
        .i* P�����������������������������������ފ            k-R�������������������������������߽j*                                                                                                                                                                                                                                    N
   N ,j
P���������������������������������������ފ.W[�͜T7DDDD����������������߆        + k����������������                          K������������������+  J    . -.JNp���������������������������������������-J          Kl�����������������������������������
MJ  
 *                                                                                                                                                                                                                              * Qi
��������������������������������������������+aC6W���W$DD&F����������������߆        + k����������������                          K������������������+  J  
 

 -Kj�����������������������������������������R          k������������������������������������� P 

                                                                                                                                                                                                                              +Ji-�����������������������������������������������kAT6�ͩ}?&&DF����������������߆        + k����������������                          K������������������+  J  
   +R�������������������������������������������k         ���������������������������������������  *                                                                                                                                                                                                                               .  kp�������������������������������������������������bA^^v���C?&&DF����������������߆        + k����������������                          K������������������+  J * ,
 
��������������������������������������������-         ���������������������������������������  *                                                                                                                                                                                                                                JJ ����������������������������������������������������,yUW���CCDF����������������߆        + k����������������                          K������������������+  J  + * ����������������������������������������������pJ         ���������������������������������������P                                                                                                                                                                                                                                  ,+������������������������������������������������������^^[���`$%&D����������������߆        + k����������������                          K������������������+  J - 
 q�����������������������������������������������J          �������������������������������������� 
                                                                                                                                                                                                                               *P �������������������������������������������������������5W����C$'F����������������߆        + k����������������                          K������������������+  J .+*-   �������������������������������������������������         Mi��������������������������������������

 
 
                                                                                                                                                                                                                             rM *l������������������������������������������������������5[[���C<'F����������������߆        + k����������������                          K������������������+  J R*-K   �������������������������������������������������        k R��������������������������������������+
 

                                                                                                                                                                                                                               . �������������������������������������������������������wT���v(H����������������߆        + k����������������                          K������������������+  J     P��������������������������������������������������R 

+ Q����������վq   ���������������������                                                                                                                                                                                                                                  J ������������������������������������������������������`[~��}8(h����������������߆        + k����������������                          K������������������+  J  
  M���������������������Ƌ�q,�l�����������������������  

, * ��������Ɋ.K+  +P�������������������                                                                                                                                                                                                                                 *  -�������������������������������������������������������8x���W2!]����������������߆        + k����������������                          K������������������+  J    M������������������߾k JM-MMi���������������������  
- , M�����הJ.QM   +Mi. ������������������                                                                                                                                                                                                                                   � ������������������������������������������������������4`���W6(H����������������߆        + k����������������                          K������������������+  J *   l�������������������Pk.    ij �������������������
   P*N* l��ߗR.P*      + i������������������                                                                                                                                                                                                                                

 JJk�������������������Ɣj,k-Q��������������������������z_���`U>>����������������߆        + k����������������                          K������������������+  J .   J������������������� J-  J  
 ii������������������-, - +M ��i, 
  *M*   KJp������������������                                                                                                                                                                                                                               -   P�����������������q  N., PP+ Q���������������������ڙ`xͨ{U=����������������߆        + k����������������                          K������������������+  J M  R�������������������  .J KR     *K������������������i  
.  . .* +
     ,i i������������������ 
  
                                                                                                                                                                                                                            KJ +P Nj������������ֽi P-  -   JN-.,����������������������vW���[=����������������߆        + k����������������                          K������������������+  J Q  +Q������������������P      ,i, *+
  ������������������q 
 
*  J.N
  + M*M��������������������                                                                                                                                                                                                                                q  P,* r����������޽i*lQiM
--
ppj.
  
����������������������W`���[>����������������߆        + k����������������                          K������������������+  J i  -P�����������������qp.    *QP , K ������������������ 
 ,. Q.*   lR*  -iiMr����������������������                                                                                                                                                                                                                                          �������ܿQ 
*                 *
��������������������G(���~`W����������������߆        + k�����������������S                        K������������������+  J -  M������������������                 �����������������   
 * . . - MP*    Q������������������������� M* 
                                                                                                                                                                                                                                     .Q������p   ,-                j��������������������g'{���[T����������������߆        + k����������������/!                        K������������������+  J -  M�����������������p                 �����������������   
 *, i    -J���������������������������� P
-  
                                                                                                                                                                                                                                    JM ����*NK*   .                  ��������������������r`���[U����������������߆        + k�����������������/                        K������������������+  J -  M�����������������N                 ������������������   
 -R  P   +p����������������������������Q*M +                                                                                                                                                                                                                                        p ��rJN PM                   �������������������߇v���v[����������������߆        + k�����������������S+                        K������������������+  J -  M�����������������-                ������������������ 
 
 .*   PMJ������������������������������ .*
                                                                                                                                                                                                                                        JpPkj J  +                 pq�������������������v{��~v����������������߆        + k�����������������/+                        K������������������+  J +  M�����������������J
                ������������������ 
    -+*R l������������������������������   * -                                                                                                                                                                                                                                        +,R J    .                 J ��������������������r`[���v����������������߆        + k�����������������"                        K������������������+  J , 
 M�����������������J                 ������������������ 
 -   -q ������������������������������� R-  +
*J                                                                                                                                                                                                                                     k *+  i .M  K
 -                Q ��������������������j'`:���x����������������߆        + k�����������������                        K������������������+  J , 
 M�����������������.                 ������������������
 
 l   JNK������������������������������
p P   --                                                                                                                                                                                                                                     lp  P-  kPN- -J                 M���������������������G(w:���|����������������߆        + k�����������������/                        K������������������+  J , 
 M�����������������J                ������������������


 
 rR 
i����������������������������� i Mk+
 -                                                                                                                                                                                                                                                     +J,   * Pi����������������������s33x�������������������߆        + k����������������׆SB-   

 M-,
P          K������������������+  J - 
 P�����������������- 

  
        ������������������ *- .
����������������������������l
                                                                                                                                                                                                                                                                     .qRr�����������������������E 7v�������������������߆        + k������������������Ar  *    M-          K������������������+  J - 
 P�����������������-     
        ������������������ -
����������������������������l. *
                                                                                                                                                                                                                                                             JN*      jjk������������������������y%%W�������������������߆        + k������������������b?,-*   *  ---P        K������������������+  J - 
 P����������������� j             ������������������  + ������������������������ֽrK  ,                                                                                                                                                                                                                                                               M     P .M��������������������������%$T~������������������߆        + k������������������b    -   P   -        K������������������+  J - 
 P�����������������,M   
           ������������������  
���������������������ֽjJM
                                                                                                                                                                                                                                                                  ,J p���������������������������1F):`������������������߆        + k�������������������mO+,
    iJ.P         K������������������+  J - 
 P������������������i  
          ������������������ 
  l�������������������R ..  
   
                                                                                                                                                                                                                                                               KpN k�����������������������������24F)V_������������������߆        + k��������������������a
  * *QJq         K������������������+  J - 
 P�������������������   
          ������������������ 
 ������������������ PM  ** -J   
                                                                                                                                                                                                                                                             M- q������������������������������z:1%D)	:_������������������߆        + k���������������������M *.  J
- ��+        K������������������+  J - 
 P�������������������-
           ������������������ *,�����������������NliR   NN 
    J                                                                                                                                                                                                                                                            j-r�������������������������������o]::%F)7Zv�����������������߆        + k����������������������p*  
�������
        K������������������+  J - 
 P�������������������J          ������������������ J.����������������RiK iR-     P*  

                                                                                                                                                                                                                                            
   

J*P  ���������������������������������q 	E	":4������������������        + k�������������������������������������M + . K������������������+  J - S�������������������                ������������������ J �����������������  +        i���J
                                                                                                                                                                                                                                               

-
*P- M���������������������������������,	J'	"1:4������������������        + k�������������������������������������.**   *K������������������+  J - S����������������֊
                ������������������ - �����������������j Mr*KQP-q�����jP--                                                                                                                                                                                                                                              
       ����������������������������������r  .. =o�����������������        + k��������������������������������������  
K������������������+  J + 
 S�����������������-                ������������������  . j����������������ʖrQkik��������� -                                                                                                                                                                                                                                                 
.*����������������������������������p+++
9Z�����������������        + k��������������������������������������. * K������������������+  J + 
 S����������������� Q                ������������������   N.���������������������������������Q,                                                                                                                                                                                                                                                
. l����������������������������������Q. E''<�����������������        + k��������������������������������������P  - K������������������+  J +  P�����������������
                 ������������������   M��������������������������������ܾ                                                                                                                                                                                                                                              
  
  -����������������������������������J  'EM<B�����������������        + k���������������������������������������- *  K������������������+  J +  P�����������������j                 ������������������ 

 *J���������������������������������p.                                                                                                                                                                                                                                            


   ����������������������������������r P
-]<'Fe&IS�����������������        + k����������������������������������������*Q  K������������������+  J )  S�����������������-                ������������������ P ,��������������������������������߽.                                                                                                                                                                                                                                            

 Pp���������������������������������* NmO,)KFe'EP�����������������        + k����������������������������������������M J K������������������+  J )  S����������������� J                ������������������ p   jQ���������������������������������i                                                                                                                                                                                                                                            +  QP�������������������������������i        e')������������������         r����������������-�����������������������.* 
K������������������M *  IPR +�����������������K.                �����������������   -
 , *��������������������������������� .* *                                                                                                                                                                                                                                      -  j-������������������������������N -        FM������������������          l����������������  ����������������������
-*-�����������������-   - )A�����������������*+                ������������������-  -+     l��������������������������������K  ,  *                                                                                                                                                                                                                                     +K����������������������������ו lR           E������������������          k���������������ߖi��������������������߅ +
�����������������*
 ,* �����������������K                ����������������֔.**   
  
 l������������������������������׽p 
.                                                                                                                                                                                                                                        iPM��������������������������ņ              MEr����������������        QQ����������������
-r��������������������M ,*�����������������rKJ

Q<�����������������Q                ����������������Ն JQ    *+  .RJ*����������������������������Օ   


                                                                                                                                                                                                                                       R������������������������ܽi
JK  . K            M   "O����������������֋         r���������������߽ X����������������֖  * �����������������q -Q,,�����������������,*                �����������������M  P   KM-J*J�����������������������޾p*P,NM  -*                                                                                                                                                                                                                                     **,����������������������޾Q,i- R              +   "]��«ycob�qq�plrK        +  lpj�q��������pjli..++\n7n�������������k
R P PQkiRjpj��������Pk M- 	<anc���o�z�r�kP-ir P                M�lq�rq���������N
 .+    
M,

 ++JQ+����������������ֿ�i ,iK+   *JJ                                                                                                                                                                                                                                     Q+ ���������������������޾qjkJ  ,J  +N
             R<m]]`���@3C\$          ,   KNK        
P
   *JX]c3��c�������sIM.K 
  *--,         i.    .G" @b8��(i** 

                  J               li      
M
JR
 ..Q..Rq����������i.
K., N,  P                                                                                                                                                                                                                                    lJ ��������������������ܔl*  JJMJ.,                �S39a}���dV @mm
GE        j M Q   ,,,,,,,,QK -MJcX8:yΓ@bb\B.EEFQP*   Q-
J 
********Q 
  jg<3@�� \]OGSj++   *                 K K *,,,,,,,,rN     jN J, * kM.  *
PN-****QPJ+****jQR  + -

 
*                                                                                                                                                                                                                                    M K�������������������*                 
*.Q
                 Cd���uTT##))&&!                                F&7`��xZ4E        - 
    
          DF3Z8Z�oM,0                                                                                                                                                                                                                                                                                                                                    K j������������������                 *  
*  
                $`���v66%DD!                                D&3:���@4$%        *
   
**          &F,34d`�b$                                                                                                                                                                                                                                                                                                                                    J �������������������K                   ,                 $$���xW[M?%"5                                %%34ZİZ:B0'         
               %F<44`��@$,                                                                                                                                                                                                                                                                                                                                     . ������������������k
l                 N     ,M                $9�͸�TT&&!                                %& 4V��:B+F         

 ,--
           %F"8V@�c7                                                                                                                                                                                                                                                                                                                                      . ������������������J+,                 K  *  P                7$x���44                                F 3Yw��Z8 '        
   +,   


        F74:�� 7+ 
"                                                                                                                                                                                                                                                                                                                                    J ������������������PM -                 

Q                   CC`���Y65>                                E93Y8��78(        
  

   M  

          FD7 34�d\9                                                                                                                                                                                                                                                                                                                                    N ������������������l.J                 
J  �J                 Z���c1++1                                <!$9 ���V:          .  +   

        PB:c�:mA  +"                                                                                                                                                                                                                                                                                                                                    M p�����������������-                 jNN��pij                aC_�����ǘp33                                ]B@ ��`:38!        .
 
  R����Ɩp*         i,bZ�y_OB ,                                                                                                                                                                                                                                                                                                                                    M ������������������M.J         ..j�����Jj+  . 
   * K]S����������z]B  ,  *                         ���`4:"         
RKi���������ӆ
RJ-K  .$$ y�4a		                                                                                                                                                                                                                                                                                                                                     -������������������� QM.
     P.Mj.��������P  --  . 
  
. p�������������BB 

 

 
                        W��`:V"        M l������������� - +   ��8@		                                                                                                                                                                                                                                                                                                                                     K
��������������������� .J+   J������������N+  - 

 N
  *-p��������������$   ,                          11%%4���TT3        Qi�������������֔ K  K ZV�y:%%		                                                                                                                                                                                                                                                                                                                                     P ����������������������Ǖ�pr�����������������   M- - M*
 KK����������������   +                          11%%W_��[[3        i ���������������݇  * Z��VX%%		                                                                                                                                                                                                                                                                                                                                     *K�������������������������������������������� MM - - ** +������������������K  -                         22&&		4d���x4        J������������������  K 7Y�yT=%%		                                                                                                                                                                                                                                                                                                                                      J�������������������������������������������� 
J     
,
+������������������+ 
 .                         22&&		4Z[��[X        N������������������* @y�:V3%%		                                                                                                                                                                                                                                                                                                                                    N PR��������������������������������������������K K 
K  *r������������������� * 
                          22DD_4U��{n        ��������������������--, 9@��4:%%%%		                                                                                                                                                                                                                                                                                                                                    l  p��������������������������������������������M  K i  �������������������� 

                          22DD`4Uv��]        ��������������������QM  YZ�`V23%%%%		                                                                                                                                                                                                                                                                                                                                    K   ��������������������������������������������-i
  
 M--��������������������,R   
                        93��}[5((FF&D��������������������)R y��VB                                                                                                                                                                                                                                                                                                                                     *+ ,.��������������������������������������������  
M  J,i ��������������������KM                             03\d��[5((FF&D��������������������.. KY�Y497                                                                                                                                                                                                                                                                                                                                     .   M ��������������������������������������������-P-   *M.��������������������P.                             	3]4��x4;!'F%F��������������������A$y�17                                                                                                                                                                                                                                                                                                                                    
*  R �������������������������������������������  +,K ��������������������J                            0	=BWw��=;!&F&D���������������������yY4""                                                                                                                                                                                                                                                                                                                                      M  J������������������������������������������� * *, *������������������   
                        G	=`V��c783(''J������������������ 9y�n7A                                                                                                                                                                                                                                                                                                                                      -+   . *�����������������������������������������  NM.,   ������������������p  .- 
                        EEZZ���V33('%J������������������b7B��89<                                                                                                                                                                                                                                                                                                                                    P. .  M 
*pl�������������������������������������q
KJ  *R  *+���������������Ֆj  NJ 
                        eM8Yd��d8: lM���������������֡B7@��\\<                                                                                                                                                                                                                                                                                                                                    p-  P  j .-���������������������������������ԕriJ.
M  i*  iQ���������������)l  MM
+
                        r'"@@@��:8!Qjr���������������B\b��c b                                                                                                                                                                                                                                                                                                                                            J
*J P����������������������������־rJM                ��������������%                                (  CZ��V8]<$?��������������OBZZ�_	                                                                                                                                                                                                                                                                                                                                             +  M  ������������������������꿅P-
                  �����������AIE                                '!!9C���411<S?a���������Ȋ<\9V��1	                                                                                                                                                                                                                                                                                                                                            
+   .*-,r������������������Ɩ� +                   a$k��������cYp(                                ''(?x��T61=AMj����ҽ�P<\:��:                                                                                                                                                                                                                                                                                                                                            
    M,   .����������ǽ�jK-,*,-                     ae%%"]4���y1]                                '$[��w62OO?# 
]<AM-+O99��:V                                                                                                                                                                                                                                                                                                                                              M.   *+ MK PK,,KP,**+--,   
KM-                b'E&&]5w���626                                '% #[͞6=5A$AR<G,SMO B�� 8                                                                                                                                                                                                                                                                                                                                            -   
-MK  *  M **            
*                FDD=;66���W26                                %
#[[��a>?$ "$ma�b Z                                                                                                                                                                                                                                                                                                                                            -.-
    
 *         

        JP.                  A%%DF5X[[���v6U                                '%%#[W�Ñ^S]A b!!NPS��3:                                                                                                                                                                                                                                                                                                                                            pR
   .NJ     JJJ..JJJNJ-
M-                    qRFFFF{v���x^U                                '%&`WU��n;oOA+ ]ggG0GG0aN<�b_3                                                                                                                                                                                                                                                                                                                                                                                                    ;;##&&>>W���V8%%                                  H!V���:4D%#6U##(:7��BG                                                                                                                                                                                                                                                                                                                                                                                                                    ;;##&&>>W���Y:%%                                  H;:_��XX&%#9$U6#(1V:�d9                                                                                                                                                                                                                                                                                                                                                                                                                    55&&>>W���wW%%                                ;V8��w` 22#!9Vy�@$'                                                                                                                                                                                                                                                                                                                                                                                                                    55&&5XVx���W%%                                @d`��`$$22#((49@��@9(                                                                                                                                                                                                                                                                                                                                                                                                                    DD5hTW���`   %%%%                                 m6��x@@"(3   "53y�@9'                                                                                                                                                                                                                                                                                                                                                                                                                    DD>gTT���v    %%%%                                T{��@7"((  8��<90                                                                                                                                                                                                                                                                                                                                                                                                                    &&HhT6|��~84%%%%                                )#!!TT��vZ1F'
4c�yA$E                                                                                                                                                                                                                                                                                                                                                                                                                    &&gHT6W���:4%%%%                                i!!TY���`F'

 X��ZB<                                                                                                                                                                                                                                                                                                                                                                                                                    (11U���[6 %'F%                                D'=1V��`62!(?.EB@�cB                                                                                                                                                                                                                                                                                                                                                                                                                     ('11W���{T %&%                                ''>:���22!!)E$9��X3                                                                                                                                                                                                                                                                                                                                                                                                                     !!''W[���T:4!%&                                " _��T64 '(<@��4                                                                                                                                                                                                                                                                                                                                                                                                                    !!''(WT���[V4"'                                "97��WX9
 M$9d�d8"                                                                                                                                                                                                                                                                                                                                                                                                                    ((##)DD>]���xW:"                                22 Ac��`V@S@��Z91!(                                                                                                                                                                                                                                                                                                                                                                                                                    ((##IDD6n}���V:                                >>AZ��}::G$$d�Y@1                                                                                                                                                                                                                                                                                                                                                                                                                    !!((##I#DDHgv���VT                                 ^^FDXz��V:!!GB��@                                                                                                                                                                                                                                                                                                                                                                                                                     !!((##))DDhH[���VT$                                ^^#FF=\��Z@;!g\�yZ 1((                                                                                                                                                                                                                                                                                                                                                                                                                    Xzϣv`CC&F&&!!                                11  a���wV84c4y�B7                                                                                                                                                                                                                                                                                                                                                                                                                    3]���`C9&f&&!!                                11  =Y��w`841@��9O                                                                                                                                                                                                                                                                                                                                                                                                                    73���vV@%E&&''                                11XT���`:bB��]                                                                                                                                                                                                                                                                                                                                                                                                                    9 3���xZ@%D&&''                                116Y��@ X��B$                                                                                                                                                                                                                                                                                                                                                                                                                     =����_V&&''                                !!=4:��y_ O�\O                                                                                                                                                                                                                                                                                                                                                                                                                    ,=|���`8&&''                                !!<:8_��CaL                                                                                                                                                                                                                                                                                                                                                                                                                    0<v���xT&&''                                <=a��n�j""                                                                                                                                                                                                                                                                                                                                                                                                                    ,""<v���}W&&''                                ]XC����"                                                                                                                                                                                                                                                                                                                                                                                                                    [u���W2^&&                                %O=A����� m]$%%%                                                                                                                                                                                                                                                                                                                                                                                                                    Uu���[6T&&                                (''% O�����݊<A+                                                                                                                                                                                                                                                                                                                                                                                                                            6Y���xW6''		                                ' ==SA�����0$7\P%E                                                                                                                                                                                                                                                                                                                                                                                                                            T^x���WU''		                                (  9=9=��j���iMO$3BnI                                                                                                                                                                                                                                                                                                                                                                                                                            >=`���UU!!22                                ;!
Xn�pAeS7B�Y:]7E                                                                                                                                                                                                                                                                                                                                                                                                                            55[���[U!!22                                (!( :c��Rt#e%,Bď\\<E                                                                                                                                                                                                                                                                                                                                                                                                                            ;(W��U((66                                (!"9��X:$A)'V:��3q                                                                                                                                                                                                                                                                                                                                                                                                                              HHT`���[((66                                >;"!Bo�cY19)jI1cby��ON                                                                                                                                                                                                                                                                                                                                                                                                     81;H���|6T&D)5;                		G0F'Y@9a��   B:��YWW$M%%%%                                                                                                                                                                                                                                                                                                                                                                    11(H���~TT&&55                		'E0'EFYb8��\    9Y:��cW39<$0%%%%                                                                                                                                                                                                                                                                                                                                                                    11(H{���TT%%;5                ,,/\8\�oa   $mB4��  9 <,                                                                                                                                                                                                                                                                                                                                                                    41(Hv���WT&%55                +NXc�bB]   <\1B2��n9\B"		%%                                                                                                                                                                                                                                                                                                                                                                      T1(;`���vT)55                  <<]9@��B\   P ]o�� B 		                                                                                                                                                                                                                                                                                                                                                                              Y1!(`��T'5;                  $<7az�7\99 N$3\9��]B9

                                                                                                                                                                                                                                                                                                                                                                            a2G_Y���['5                    \9BX��n9<P ).9nXn��3                                                                                                                                                                                                                                                                                                                                                                          c6gZ:���[E5                    \b\y�z\B9$$OIP)   aBa��X                                                                                                                                                                                                                                                                                                                                                          G,EE                6U +$���~Y %%=                 M. B$\9c�cZ9y�n39:,, .                                                                                                                                                                                                                                                                                                                                                        *E<P)P0                UT
  x���@:%%>                Q   N az�Xc 9\��99B,<<                                                                                                                                                                                                                                                                                                                                                          	 ,<0L" /L,,0/,                X6+ *U���VZ&D                 *N/A<��\9X��a:Y8=9O0                                                                                                                                                                                                                                                                                                                                                          
 "<"] ]RN                U2- **U���_ZFD                
PN$B��aB9"$9 7Bc��3@\ ,                                                                                                                                                                                                                                                                                                                                                          -
  <O]ay�4n�οOO9<"""                U2#%%U{��}WfD                "OO]��O$O   
!0 B83��c8X9=9                                                                                                                                                                                                                                                                                                                                                       z�y�����]"A9A<                U2)WU���TfD9                Oa$�oo<B  **
!@\aybX39                                                                                                                                                                                                                                                                                                                                                    <$A=��a44��������o                  ^2#%&U6���[fDB                5=]��"O<"!eI' ",]39:\��V@:\                                                                                                                                                                                                                                                                                                                                                    $n��\8B:44c�����a]���b  99                ^2##DD66���vfFB                3O��<=p],!OeI)) Obb���89                                                                                                                                                                                                                                                                                                                        %%	 NA1X41c��B %%5�����]"o��y86Y411883<O'%FF%&22|���V8#'')
 $VY8��                                                ]a��@B                                                                                                                                                                                                                                                                                                        D'  A9bb>1y��Tb 5d�ď"<A99���21113B<G"%'%&22u���Z8G0'''F%'9@Z2��a                                                1]X��7@B<G                                                                                                                                                                                                                                                                                                            $$A\ b��z1VB	34��VY<aA$$a��z48B="OGM%%  [���`WM)  V�o9N                                                =anĈ77<<"                                                                                                                                                                                                                                                                                                          ) ,<<BB��o\:BV134��4:"\\ ���\ <L%%[����V#<<0,'97@b�4a <                                                =]@ ��B 9=<N                                                                                                                                                                                                                                                                                                              <AA$O$\��<"093  $9	":��Y8,<$?95]���9]]11T`�͞4$<AbBn� BA,]                                                <OB] z�aX\:4                                                                                                                                                                                                                                                                                                              $O<��<9]BOB\7 0X��22]"0/A]$<=B93z��]<<On11[:���`"$""",nB��9 9A<M                                                 <=9=\7 48:\                                                                                                                                                                                                                                                                                                          9B9Bn��nO]O"  <b)$3c��V2 *G]<A"=���=Xb:62_9���y=$" 9 9a\��aOO""e%                                                "GLA]9n3��c1ZV                                                                                                                                                                                                                                                                                                          Cb9B��o�]<<7 ""JKA)$:zЂYV\XjR+O<"97 �aXy��o866@9`wVWo���ˏ]r$n�o9B9m -*M                                                iOB 9XcY��1Y                                                                                                                                                                                                                                                                                                    N . !RiC��o9\AV��[:4='*    Y���^,A$7@:��������9a\a�a99                                                9=X1V��Vn9LM<                                                                                                                                                                                                                                                                                                     +-
M!!]<B��\B% BV��W84<'*  14z��z,L-?a�����������7z�o                                                8@X14��oXB 0NEEi]"                                                                                                                                                                                                                                                                                                       
<,"a���B O 9'  7XW��V<%'7983]=���A$m�����������䏙]9""                                                  <3OB8:Z��9="E���p i                                                                                                                                                                                                                                                                                                    	   OmOr��B 9  )  :X[��V3(%%388XX1<z��q$��������������3=9]NL                                                  "37B:3B��ojLNp������,                                                                                                                                                                                                                                                                                                      +M<Oz��3O<O!0@Vv��@ %%26==r!��������������n=GE                                                  $$mX4\�]�������l                                                                                                                                                                                                                                                                                                      Mi���o�7\33<<<!"00@V��@3'!,<NS336:>>;O��������������O(S                                                  'O$4X]�������ݑM                                                                                                                                                                                                                                                                                                    I)+Q�����=B8SGG0		G:T��cC"F%%ME''* 3^UUU]!���������������m"R0%%                                                %%F%  *1X9n���������                                                                                                                                                                                                                                                                                                    l).E/�����n48gQGEGG(:T��b9F%%RMGE''+KB32662HO���������������],0EIF                                                %%eEFE*   y8]���������Q                                                                                                                                                                                                                                                                                                    EI)�����@\,                 %;H8W��
                                      , ��������������M,  
                                                                                 --q�������J                                                                                                                                                                                                                                                                                                    )I����  
E                %;G:[��
                                       i��������������-  
                                                                                 -*  
*P�������ij                                                                                                                                                                                                                                                                                                    $%��oa\%F                !!'5;:`��
                                      Q
 ������������q                                                                                    J*  K*N�����Q.P                                                                                                                                                                                                                                                                                                    <),nbX%E                !!E""Vw�}
                                      ,QMJ����������                                                                                       
  J- ., M 
                                                                                                                                                                                                                                                                                                     OEE"<�o1Y K                !!NV�v
                                      * , ��������i .  

                                                                                       
* M, J,                                                                                                                                                                                                                                                                                                      O<S��1Y\9'                !!SV��v
                                         QM����K*Q  

                                                                                   *  ,J   -
  *K,                                                                                                                                                                                                                                                                                                    ](']��T2\]                RV��v
                                         - M.J*jk
-                                                                                    P *N   
   *.                                                                                                                                                                                                                                                                                                    ]=<O��{T4S                QV��x
                                      l. 

  qK
  *MP                                                                                     PK 
*   lMM -                                                                                                                                                                                                                                                                                                       Y��W11S"                9@`��V                                                                                                                                                                                                                                                                                                                                                                                                                                                                    Yy�6X1]                $ @w�w:                                                                                                                                                                                                                                                                                                                                                                                                                                                                    :Z�`Y1<                 '%$@@��`6                                                                                                                                                                                                                                                                                                                                                                                                                                                                    2W��VV<                '%9@9��T4                                                                                                                                                                                                                                                                                                                                                                                                                                                                    4Yw�Y@A                '&C$7��24                                                                                                                                                                                                                                                                                                                                                                                                                                                                    VVV��37                '&C$C��24                                                                                                                                                                                                                                                                                                                                                                                                                                                                    		Z3:��8A                D'C7_��22                                                                                                                                                                                                                                                                                                                                                                                                                                                                    		Z6�ZO                D'C7@d�41                                                                                                                                                                                                                                                                                                                                                                                                                                                                        < a��Z2	 %% V�c8                                                                                                                                                                                                                                                                                                                                                                                                                                                                        "B��WT
%% V��c8                                                                                                                                                                                                                                                                                                                                                                                                                                                                        "y�`Z%%:V��Y7                                                                                                                                                                                                                                                                                                                                                                                                                                                                        "Y��Z!%%:V��Z                                                                                                                                                                                                                                                                                                                                                                                                                                                                          :��Y 38ZY                                                                                                                                                                                                                                                                                                                                                                                                                                                                        98b�y"81c_                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ,<7��73:1�cZ                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ,$7��73V1��Y@                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ,+<37@�cy\O1Y��@B                                                                                                                                                                                                                                                                                                                                                                                                                                                                     /$ 97��c\A1Y��@B                                                                                                                                                                                                                                                                                                                                                                                                                                                                     G"9n�cV130 2YÎ79 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                    E$9��1402c� 9                                                                                                                                                                                                                                                                                                                                                                                                                                                                     *��1:-33:w�w                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ){�VV+33W�w                                                                                                                                                                                                                                                                                                                                                                                                                                                                    E "w��Z933Y��w)                                                                                                                                                                                                                                                                                                                                                                                                                                                                    E) <{��_X33c��w)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ��`YT=%%	'(('3d��_7(;                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     Y�Y:8%%	(('3d��_7(H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    3��Y:14%%	((!3�}C (H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    33_�wT11%%	(!8��_C  (H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     @1��6:%	!! 9��CC ';                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    994y�:\%	!!39��CC7'(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    O@:�yY1	3:C97(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    b@1��V1	7@āC77(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    B@c�Z: 

<Zc�y@7B0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    B9Z��8  	5 @��d97<(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    936��:7!!3:@��@9 "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    E34y�c9 <@8��79                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     %eVW��7 !O!9@�� 9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     %IY:��8 "](37Z��9 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     IDV8w�b@(g;9 9d��@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     e&"48`��Yg;= 9���X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ((+@��`Z4OF&<$6[��V:                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ($3c�wWV<f&<$6[��V:                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    !$8��TV9I%796W��V8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    $7 ��V2  F%' 76W��:4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    8 c�w293%E7T[��:4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    !7 _��6B FM7Tw�:4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    0
   cy�cB0P 8W��{8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    <   9y1�{9/P 8[��{8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    1b��@8OS`��W		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    1Yy�XXBN1`��W		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    1:V�yV9911wV		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ::��8B714w�wT		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    %%:6y�Y@B46�`:                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    %%:92c��:X46��Y:                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    %%=2Y�Z \48��Y:                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    %%\VV`�c \44��Y:                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    +6��6^66cĉ1]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    + 2��W666c�y2]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    *994X�w26T��y4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    9V2��226��X1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      :1��\��9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      11Y�y:=��]9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    14��B S<$+                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      M::18a9<OA<$]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ��, J                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    A����K
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �����R                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �����NP                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      i����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    GGg,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    kS!R,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              BM�      �   |                    �  �            �  �  �      �BGRs                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 H�H�F�$N�"L�%O�"N�I�H�"L�'Q�%O�$O�"L�&P�"N�	*T�
+U�(R�'Q�"L�!L�H�&P�'Q�&P�'P�!L�J�"P� ! ])4y�	6{�5y�B��@��A��G��
8}�5z�?��E��B��B��?��D��C��I��J��J��F��?��>��
9}�B��G��F��C��>��
:~�@��/p; %g/
:��
:�>��I��F��G��J��
;��	8�B��J��E��D��C��H��A��P��R��P��J��E��?��=��I��K��K��K��C��>��E��7zI (n3@��=��C��O��L��I��G��>��
;��F��K��G��H��F��M��E��U��N��T��O��G��C��B��N��P��N��L��H��C��I��A�N2u=E��A��E��U��Q��Q��P��C��=��L��R��K��M��J��S��S��X��R��V��S��J��F��E��P��T��P��O��K��G��L��@�O4y?H��E��K�� Y��U��S��W��I��E��Q��X��T��Q��O��W��Y��#Z�� Y�� Z��Y��P��L��G��U��X��W��T��P��K��Q��M�O
>�JN��O��P��&_��!Z��$]��$^��M��L��U��&_��!Z��T��S��![��X��)a��(a��&`��%_��U��P��N��!Z��"\��&`��'`��"Y��M��W��S�OC�OT��W�� W��-f��)c��*c��)b��S��P��#[��+d��$]�� Y��![��(a��W��/h��/h��,f��+e��X��W��R��'`��(b��1j��-f��)a��U��"[�� Z�OK�X X��!Y��%\��1j��1j��-f��,e��W��S��&^��0i��'`��"[��$]��,e��R��3l��3l��0j��-g��#]��"Z��T��/h��.h��4m��1j��,e�� X��&_�� Z�ON�^"Y��%\��)`��-f��1j��/i��0i��#Z�� V��,c��2k��)a��$\��'`��.g��*b��6o��4n��5n��1k��*c��$[��#[��3l��2l��6o��4m��/g��$Z��)b��K�U"W�i%\��'^��*c��-f��,d��3l��5n��&]��#Y��.f��5n��.f��)a��+d��0i��2l��8q��2j��6o��8q��3l��'^��(`��7p��5n��:s��7p��0h��$[��*c��C�^"[�o(]��+a��-f��0i��0i��6p��9q��)_��'\��3j��;t��4m��-e��/g��1k��3m��8q��5n��9r��;u��7p��,d��*b��8q��6o��<u��:s��5m��(^��-e��H�i"X�|,b��,c��/g��4m��0h��9r��:s��-d��*`��7n��>w��7p��1i��1j��4m��6n��;s��7p��;u��?x��<u��0h��.e��9r��8q��:s��>w��7p��,b��1i��M�v(^��/f��1h��4l��8q��3k��=u��>v��0g��/e��:r��Az��9q��5n��5n��7p��7p��@x��?x��?x��C|��?x��3k��1h��=v��=v��@y��Az��9p��.c��0f��"V��*`��2i��5k��7p��:s��5m��>w��>w��1g��1g��=t��E~��?x��8r��9r��:r��9r��C{��?w��B{��F��C|��9r��6o��?x��@y��@y��C|��;s��3i��4k��#V��/d��4k��7n��9r��;s��9p��@y��@y��4j��1f��?w��E~��D}��=w��=v��=v��;t��D{��D}��C|��G���F~��9r��8q��>w��C|��B{��F��@x��4k��8o��'Y��0f��5k��8n��;s��>v��<t��E}��B{��7n��4i��D|��H���F��A{��@y��>v��<t��G��F��E~��H���G���;t��;s��?w��C|��C|��H���C{��7n��>v��,a��4j��6l��:p��<u��>v��=t��D}��Az��9o��5i��F|��I���I���B|��Az��Bz��:r��G��I���M���J���G���<t��<t��B{��G��G���J���F~��9o��<t��0d��6l��8n��;r��=u��<t��=t��C|��Bz��8n��4h��F~��G���F~��B{��B{��Bz��8n��J���K���O���K���H���>v��<s��F��L���I���L���I���<s��;r��5j��K��bBu��=q��?s��?u��?t��E{��Bx��=q��9j��F{��H��G}��F}��D{��Dy��?t��M���O���O���J���H}��@v��?t��H~��L���I���M���J��>s��J���M��i    /v+D��>��H��M��M��O��H��>��C��Q��J��L��I��N��J��V��W��T��P��H��G��G��M��Q��R��O��C��N��=�            <t�;S��'`��)c��&`��&`�� Y��Q�� W��)c��#^��'a��G��NY��?L��?a��?a��?]��?Y��?P��?L��?P��?Y��?Y��?]��?Y��?L��?W��                    )_��8q��=v��8r��7q��0i��)^��0h��9s��2k��1k��                                                                                    F|�^T�̿Y�пV�οT�ͿM�ȿH}¿L�ƿX�пS�ͻS��@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              BM�      �   |                    �  �            �  �  �      �BGRs                                                                                                                                                                                                                                                                                                                                      111R111�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�111�111R       $$$222�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�222�$$$333�333�333�222�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�222�333�333�333�222�333�222�                                                                                                      222�333�222�222�333�222u                                                                                                        222u333�222�333�333�222u                                                                                                        222u333�333�333�333�222u                                                                                                        222u333�333�333�333�222u                                                                                                        222u333�333�333�333�222u                                                                                                        222u333�333�333�333�222u        ///+222�333�333�+++                ...333�333�333�333�333�333�333�222�333                    222u333�333�333�333�222u            3337333�333�333�+++            ...,333�333�333�333�333�333�333�333�111S                    222u333�333�333�333�222u                3337333�333�333�+++            222`222�222�222�222�222�222�111q                       222u333�333�333�333�222u                    3337333�333�333�+++                                                                222u333�333�333�333�222u                        222�333�333�222�                                                                222u333�333�333�333�222u                    222e222�333�222�$$$                                                                222u333�333�333�333�222u                222e222�333�222�$$$                                                                    222u333�333�333�333�222u            222e222�333�222�$$$                                                                        222u333�333�333�333�222u        ///+111�222�333�$$$                                                                            222u333�333�333�333�222u                                                                                                        222u333�333�333�333�222u                                                                                                        222u333�333�333�333�222u                                                                                                        222u333�333�333�333�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�222�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�222�222�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�222�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�$$$222�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�333�222�$$$       111R222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�222�111R                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             BM�      �   |                    �  �            �  �  �      �BGRs                                                                                                                                                                                                #&&&&&&&&&&&&&&&&#                                  YY]G�������ʽ��ώ�㽽�㽽�㽽�㽽�㽽�㽽�㽽�㽽�㽽�㽽�㽽�㽽�㽽�㽽�Ḹ�ʪ���[[[F                          #������������������������������������������������������������������������������������������������#                  ��������������������������������������������������������������������������������������������������������           
���`�����������������������������������������������������������������������������������������������������������`
        ����������������������������������������������������������������������������������������������������������������       PPP)����������������������������������������������������������������������������������������������������������������PPP)      ���H�������������������������������������������������������������������������������������������������������������������H      ���K�������������������������������������������������������������������������������������������������������������������K      ���I�������������������������������������������������������������������������������������������������������������������I      ���G�������������������������������������������������������������������������������������������������������������������H      ���H�������������������������������������������������������������������������������������������������������������������H      ���I�������������������������������������������������������������������������������������������������������������������I      ���G�������������������������������������������������������������������������������������������������������������������H      ���I�������������������������������������������������������������������������������������������������������������������I      ���G�������������������������������������������������������������������������������������������������������������������H      ���G�������������������������������������������������������������������������������������������������������������������H      ���I�������������������������������������������������������������������������������������������������������������������I      ���G�������������������������������������������������������������������������������������������������������������������H      ���H�������������������������������������������������������������������������������������������������������������������H      ���M�������������������������������������������������������������������������������������������������������������������M      C<9L�|w������|w������|w������|w������|w������|w������|w������|w������|w������|w������|w������|w������|w������|w�����C<9L      2.+GB:3�C;4�B:3�C;4�B:3�C;4�B:3�C;4�B:3�C;4�B:3�C;4�B:3�C;4�B:3�C;4�B:3�C;4�B:3�C;4�B:3�C;4�B:3�C;4�B:3�C;4�B:3�C;4�5.+G      1,(9C;4�B:3�B:3�B:3�B:3�ZSM�����������������������}�NF@�������������������������ke_������}x�f_Z�B:3�B:3�B:3�B:3�C;4�0+':      D<5�D<5�B:3�B:3�B:3�d]W�d^X�PHB���������oic���������������������a[U�����������������\UO�D<5�B:3�B:3�B:3�D<5�D<5�       A93�F>7�E=6�B:3�B:3�B:3��}y�����zto�mga�|wr�tni�upk�rlg���}�����������������������~�B:3�B:3�B:3�B:3�E=6�F>7�A93�           ,,'4F>7�G?8�G?8�F>7�D<5�����pid�����D<5�D<5�D<5�D<5�D<5�D<5���~�����D<5�TLF�����g`[�D<5�D<5�F>7�G?8�G?8�F>7�1,'4               930YG?9�H@:�H@:�H@:�PIC�ysn�WPJ�H@:�H@:�H@:�H@:�H@:�H@:�KD=�mga�H@:�H@:�����jd^�H@:�H@:�H@:�H@:�G?9�930Y                   73,EF@9�IB;�IB;�IB;�IB;�IB;�IB;�IB;�IB;�IB;�IB;�IB;�IB;�IB;�IB;�IB;�IB;�IB;�IB;�IB;�IB;�F@9�73,E                          85.HC=7�E>7�E>8�E>8�E>8�E>8�E>8�E>8�E>8�E>8�E>8�E>8�E>8�E>8�E>8�E>8�E>7�C=7�85.H                                         

                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                BM�      �   |                    �  �            �  �  �      �BGRs                                                                                      T   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   U                                          �   l   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   k   �                                      @   �                                                                                   �   @                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �                                                           L   y   {   {   {   {   �   B                                   B   �                                                       �   �   �   �   �   �   �   �   8                                   B   �                                                      �   G                  �   �                                       B   �                                                   	   �   %              �   �                                          B   �                                                   	   �   %          �   �                                              B   �                                                   	   �   %       �   �                                                  B   �                                                   	   �   %   a   �   1                                                   @   �                                                   	   �   g   �   M                                                          �   l   /   /   /   /   /   /   /   /   /   /   /   7   �   �   n                                                               T   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  BM�      �   |                    �  �            �  �  �      �BGRs                                                                                      T   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   U                                          �   l   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   k   �                                      @   �                                                                                   �   @                                   B   �                                                                                   �   B                                   B   �           .   B   B   B   B   B   B   B   B   B   B   B   B   B   B   .           �   B                                   B   �           �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �           �   B                                   B   �                                                                                   �   B                                   B   �                                                                                   �   B                                   B   �           ~   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ~           �   B                                   B   �           V   z   z   z   z   z   z   z   z   z   z   z   z   z   z   V           �   B                                   B   �                                                                                   �   B                                   B   �              %   %   %   %   %   %   %   %   %   %   %   %   %   %              �   B                                   B   �           �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �           �   B                                   B   �              	   	   	   	   	   	   	   	   	   	   	   	   	   	              �   B                                   B   �                                                                                   �   B                                   B   �           j   �   �   �   �   �   �   �   �   �   �   �   �   �   �   j           �   B                                   B   �           j   �   �   �   �   �   �   �   �   �   �   �   �   �   �   j           �   B                                   B   �                                                                                   �   B                                   B   �              	   	   	   	   	   	   	   	   	   	   	   	   	   	              �   B                                   B   �           �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �           �   B                                   B   �              %   %   %   %   %   %   %   %   %   %   %   %   %   %              �   B                                   B   �                                                                                   �   B                                   B   �           V   {   {   {   {   {   {   {   H               L   y   {   {   {   {   �   B                                   B   �           }   �   �   �   �   �   �   �   j           �   �   �   �   �   �   �   �   8                                   B   �                                                      �   G                  �   �                                       B   �                                                   	   �   %              �   �                                          B   �           �   �   �   �   �   �   �   �   �       	   �   %          �   �                                              B   �           .   B   B   B   B   B   B   B   '       	   �   %       �   �                                                  B   �                                                   	   �   %   a   �   1                                                   @   �                                                   	   �   g   �   M                                                          �   l   /   /   /   /   /   /   /   /   /   /   /   7   �   �   n                                                               T   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ELF          >       �   @       8t         @ 8  @  
                 �      �    �       �                    �       �  �    �  �   x        0                            �      �                          Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��  ���_ cole _          �      �            @ �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           I��H�p �   L�H�P �   H�H� �  �   L�H��  �   L�#H��  �   L�+�   �����H��H��H��H��L�������UH��AWSH��@��H�����I���      L�H�}�H�u�H�U�H�M�L�E�L�M�H���������H�H�U�H�H�     H�E�H�H�E�H��     H�H��     H�H� H��H�      H�H��     H�H��H��     H�H��     H�H�@H��H��     H�H�E�H��     H�H�E�H��     H�H�E�H��     H�H�     H�H��H��     H�I�߸    H��G������H���H��     H�    H���������H�H� H��H��     H�H���������H�H� H��H���������H�H� H�։�I��H��������H��ЉE�E��I��H�f�������H��АH��@[A_]���UH��AWSH�� ��H�����I��      Lۉ}�H�u�H��������H�fHn�I��H�h�������H����E�H� �������H�fHn�I��H�h�������H����M�H��������H�<I�߸   H�r�������H��Ҹ    H�� [A_]���UH��AWSH����H�����I�`�      Lۉ}�H�u�H�E�� ��H�E��@9�sH�E��P#H�E��@9�r"H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@��u)H���������H�H��E�H�։�H��������H���H�E�H�PH�E��@#��H�H�E�H�PH�E�H�@�U�H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  H�E��@��u0H���������H�H� H��t�E�����I��H�Df������H��ЋE�H��[A_]���UH��H����H�����I�	�      L�H�}��E�    H�E�@��u]H�E�@'�PH�E�P'��H�E�P#H�E�@'9�r�H�E�H�PH�E�@'��H��H�H�E�H�PH�E�H�@� ���E��   H�E�@��tH�E�@��uiH�E�@#��u������ZH�E�P'H�E�@#9�r������AH�E�H�PH�E�@'��H�H�E�H�PH�E�H�@� ���E�H�E�@'�PH�E�P'�E�����UH��H����H�����I���      L�H���������H�H� H�E��E�    H�E��@��uWH�E��P#H�E��@'9�w�    �AH�E�H�PH�E��@'��H�H�E�H�PH�E�H�@� ���E�H�E��@'�PH�E��P'�E�����UH��H����H�����I�C�      L�H���������H�H� H�E��E�    H�E��@��uXH�E��@'�PH�E��P'��H�E��P#H�E��@'9�r�H�E�H�PH�E��@'��H��H�H�E�H�PH�E�H�@� ���E��E�����UH��AWH��(��H�����I���      L�H�}�H�u�H�U����u�    �(H�M�H�U�H��H��I��H�1.������H���H�E�H�E�H��(A_]���UH��AWSH�� ��H�����I�'�      L�H�}�H�}� u
������   H�}� tH�E؋@����tH�E��@"<t������zH�E؋@%�   ��u�    �cH�E؋@#H�U؋J�    ��E�H�E؋@��@��u�U�H�E؉�H��I��H��8������H���H�E�H��I��H�u5������H��ЉE�E�H�� [A_]���UH��AWSH����H�����I�@�      L�H�}�H�}� u������0H�E�H��H��������H���H�E�H��I��H��6������H���H��[A_]���UH��AWSH�� ��H�����I���      Lۉ}�H�u�H�}� u
�������  H�EЋ@��u
�    �  H�EЋ@��tH�EЋ@��tH�EЋ@��u!H�UЋE�H�։�H��������H����y  H�EЋ@����unH�EЋP#H�EЋ�+  9�wYH�EЋ�+  ��tKH�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��E�U�H�EЉ�H��I��H��7������H����H�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U܈H�E�� ��H�EЋ@��9�r3H�EЋ@����H�EЉPH�E�f�   H�E�H��H��������H���H�EЋ@#�PH�EЉP#H�EЋP#H�EЋ�+  9�vH�EЋ�+  �PH�EЉ�+  H�EЋ@���H�EЉP�    H�� [A_]���UH��AWH��(��H�����I���      L�H�}�H�}� u
������  H�E؋@��u
�    �v  H�E؋@��tH�E؋@��tH�E؋@��u"H�E�H��H��������H��ЉE�E��0  H�E؋P#H�E؋�+  9�r
������  H�E؋@����ulH�E؋P#H�E؋�+  9�wWH�E؋�+  ��tIH�E؋@����H�E؉PH�E؋@#H�U؋r�    ���E�U�H�E؉�H��I��H��7������H���H�E؋@#H�U؋J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@� ���E�H�E�� ��H�E؋@��9�rH�E؋@����H�E؉PH�E�f�   H�E؋@#�PH�E؉P#�E�H��(A_]���UH��SH��H��H�����I���      L�H�}ȉuĉU�H�M�H�}� u�    �y�E�    H�E�H�E��E�    �FH�E�H��H�?������H��ЉE؃}��u�E�    �u��4H�E�H�PH�U��U؈�E��E��E��E��E�9�w��E�    �u�H��H[]���UH��SH��H��H�����I�$�      L�H�}ȉuĉU�H�M�H�}� u�    �l�E�    H�E�H�E��E�    �9H�E�H�PH�U�� ���E�H�U��E�H�։�H�#������H��ЃE��E��E��E��E�9�w��E�    �u�H��H[]���UH��H����H�����I�q�      L�H�}�H�u��U�}�tZ�}�|�}� t�}�t�nH�E���H�E��P#H�E���H�E��P'�RH�E��@#H�U��H�E��P#H�E��@'H�U��H�E��P'�(H�E���+  H�U�)Љ�H�E��P#H�E��P#H�E��P'�H�E��@#H�U��J�    ��Љ�H�E�f��    ����UH��H����H�����I���      L�H�}�H�}� u�    �	H�E��@#������UH��H����H�����I�R�      L�H�}�H�}� t7H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@����H�E��P������UH��H��(��H�����I���      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H��(��H�����I���      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H����H�����I�?�      L�H�}��E�_   �(�E�Hc�H�E�H�� < u�E�Hc�H�E�H��  �m��}� y����    ����UH��H����H�����I���      L�H�}�H�E�H�E�H�E�H�E��H�E�� </uH�E�H��H�E�H�E�H�E�� ��u�H�E�����UH��H��0  ��H�����I�l�      L�H������H������H������H�E�H������H�E�H������H�E��E�    �?H�E�� ��u�E�Hc�H�E�H��  �H�E�H�PH�U��U�Hc�H�U�H�� ��E��}�_~��E�    �-H�E�H�PH�U��H�E�H�PH�U�� 8�t�   ��E��}�_~͸    ����UH��SH�� ��H�����I���      L�H�}�H�u�H�E؋PH�E؋@ЉE�E�H�U����H�@     H�H�¾   H�������H��ЉE�}� t
�������   �E�    ��   �E�%�  ��H�@     ��H؋���uf�E�%�  ��H�@     ��H��������E�H�U����H�@     H�H�¾   H�`������H��ЉE�}� t������r�E��m�E�%�  =�  uE�E��E�H�U����H�@     H�H�¾   H�������H��ЉE�}� t�������E�H�E؋@$9E����������H�� []���UH��H����H�����I���      L؉}��u�H�U�H�M�    ����UH��AWSH��0��H�����I���      Lۉ}�H�u�H�U�H�EȋPH�Eȋ@ЉE�H�Eȋ@ �E܉E�ЉE�   �    H�@     H�<I��H��t������H����E�    �B�U�E�Љ�H�EЋ ��H�@     H��   H�`������H��ЉE��}� u�E�H�EȋP �E�9�w���H��0[A_]���UH��H����H�����I���      L�H�}�H�u�H�U��R��H�U����H�U�H��H��   I�������J� ������UH��AWSH��`��H�����I�{�      L�H�}�H�u�H�U�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H�'�������H���H�E�H�E�H�E�H�E�H��I��H��U������H��ЉE�H�E��@,�E��9  H�E�H�E��H�E�� </uH�E��  H�E��H�E�H�E�� ��u׋U�H�E��@ H�M��	��H�M���H�������H��ЉE؃}� t#H�E�H��I��H�ö������H��и    ��   �E�    �f�E���Hc�H�E�H�H�E�H�E��@a��t5H�E��@b����@��t#H�E�H�U�H��H��H�� ������H��ЉE���E������}� t�E��}�?~����}� u+�}�?%H�EЋ@k�E�H�E��@ �E؉E�ЉE�m��	�E�    �
�}� �����H�E�H��I��H�ö������H��ЋE�H��`[A_]���UH��AWSH��P��H�����I�f�      L�H�}�H�u�H�U��M�L�E�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H�'�������H���H�E�H�Eغ    �    H��I��H��t������H��ЋU�H�E��@ H�M��	��H�M؉�H�������H��ЉE�}� t#H�E�H��I��H�ö������H��и������   �E�    �T�E���Hc�H�E�H�H�E�H�E��@a��t#H�E�H�U�H��H��H�� ������H��ЉE���E������}� t�E��}�?~����}� u:�}�?4�E���Hc�H�E�H�H�EȺ�   H��H��I��H�1t������H�����E�����H�E�H��I��H�ö������H��ЋE�H��P[A_]���UH��AWSH��P��H�����I���      L�H�}�H�u�H�U�H�E���C  ��u
������	  H�E���C  ��@v/H�(�������H�<I�߸    H�r�������H��Ҹ������  H�E��PH�E��@ЉE�H�E���?  H�E��@ �ЋE�ЉE�    I��H�'�������H���H�E�H�Eغ    �    H��I��H��t������H��ЋU�H�E��@ H�M��	��H�M؉�H�������H��ЉEԃ}� t!H�E�H��I��H�ö������H��ЋE��  H�E���C  ��H��H��H�E�H�H�E�H�EȺ`   �    H��I��H��t������H���H�E�H��+H��H� ������H���H��H�E�H��H��I��H�:w������H����E�    �"H�UȋE�H����uH�UȋE�H�� �E��}�_~�H�E��@` H�E���+  H�EȉPo�U�H�E��@ H�M��	��H�M؉�H�`������H��ЉE�H�E�H��I��H�ö������H��ЋE�H��P[A_]���UH��AWSH��`��H�����I�?�      L�H�}�H�u�H�U��S  I��H�'�������H���H�E�H�EкS  �    H��I��H��t������H���H�E��PH�E��@ ��H�EЉP�    I��H�'�������H���H�U�H�BH�E��PoH�EЉ�+  H�E��PH�EЉ�/  H�E��P H�EЉ�3  H�E��H�EЉ�G  �    I��H�'�������H���H�U�H��K  H�E�H��K  �    �    H��I��H��t������H���H�E��@k�E�    I��H�'�������H���H�E��E������E�    �E�    ��  �   I��H�'�������H���H�U�H��K  �M�Hc�H��H�H�H�E�H��K  �U�Hc�H��H�H� H�E�H�E��   �    H��I��H��t������H����E�    �<  H�E��@ �E��H�E��@�H�E��P�E�H�H�4�    H�E�H�ʉH�EЋ�;  �PH�EЉ�;  �E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E�;E�ts�E�H�U����H�U�H��H�¾   H�������H��ЉE��}� t:H�E�H��I��H�ö������H���H�E�H��H��6������H��и    �   �E��E�H�E��@�����E�    ��U�E�H��    H�E�HЋ �E�}��u	�E�������E��}��  ������}��t�E��}��  � �����H�E�H��I��H�ö������H���H�E�H��`[A_]���UH��AWSH��p  ��H�����I���      L�H������H�������   I��H�'�������H���H�E�H�E�H�E�H�E�H   H�E�H������H�E�H��H��I��H�fS������H���H�U�H�E�H��H��I��H�V������H��п�   I��H�'�������H���H�      H�H�      H���   �    H��I��H��t������H��п   I��H�'�������H���H�E�H�EȺ   �    H��I��H��t������H���H�E�H�E�H�E��   �    H��I��H��t������H����E�    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ ���    Hǅ���    Hǅ���    Hǅ���    Hǅ ���    Hǅ(���    Hǅ0���    Hǅ8���    Hǅ@���    HǅH���    HǅP���    HǅX���    Hǅ`���    Hǅh���    Hǅp���    Hǅx���    H�E�    H�E�    H������H������H��H��I��H�:w������H���������<wt������<au�E�   H�E��@   H�E��     H�U�H�E�H��H��H�$������H��ЉE�}� t_H�      H�H��I��H�ö������H���H�E�H��I��H�ö������H���H�E�H��I��H�ö������H��и    �  H�E�H�U�H�M�H�E�H��H��H�v$������H��ЉE��}� u_H�      H�H��I��H�ö������H���H�E�H��I��H�ö������H���H�E�H��I��H�ö������H��и    �  H�EȋU��P,H�      H�H�M�H�U�H�u�I�ȹ    H��H��&������H��ЉE�}����   �}� tqH�      H�H������H�U�H�u�A�    H��H�F=������H���H�      H�H������H�U�H�u�I�ȹ    H��H��&������H��ЉE�}� ��   H�      H�H��I��H�ö������H���H�E�H��I��H�ö������H���H�E�H��I��H�ö������H��и    ��  �}� t_H�E�H��I��H�ö������H���H�      H�H��I��H�ö������H���H�E�H��I��H�ö������H��и    �r  H�      H�H�U�H�M�H��H��H��*������H���H�E�H�}� ��   H�      H�H��H�E�H��+�`   H��H��I��H�1t������H���H�E�H��+H��H��������H���������<wt������<+t������<au
H�E��@"�H�E��@"H�E��@   H�EȋP,H�E���?  H�      H��PsH�E���C  ������<auH�      H��PoH�E��P#H�E�H��I��H�ö������H���H�      H�H��I��H�ö������H���H�E�H��I��H�ö������H���H�E�H��p  [A_]���UH��AWSH��@��H�����I�|�      L�H�}��   I��H�'�������H���H�E�H�E�   �    H��I��H��t������H���H�E�H�E�H�E�   �    H��I��H��t������H���H�E��@   H�E��     H�U�H�E�H��H��H�$������H��ЉE܃}� t H�E�H��I��H�ö������H��и�����AH�U�H�M�H�E�H��H��H�U(������H��ЉE�H�E�H��I��H�ö������H��ЋE�H��@[A_]���UH��AWSH�� ��H�����I�B�      L�H�}�H�E�H�@H��I��H�ö������H����E�    �TH�E�H��K  �U�Hc�H��H�H� H��t?H�E�H��K  �U�Hc�H��H�H� H��I��H�ö������H��ЃE��}��  ~���H�E�H��K  H��I��H�ö������H���H�E�H��I��H�ö������H���H�E�    �    H�� [A_]���UH��H�� ��L�����I�E�      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H�������I� ������UH��H�� ��L�����I�q�      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H�`������I� ������UH��AWSH��   ��H�����I���      L�H��x���H��p�����l����   I��H�'�������H���H�E�H�E�H�E�H�E�H   H�E�H��x���H�E�H��H��I��H�fS������H���H�U�H�E�H��H��I��H�V������H��п   I��H�'�������H���H�E�H�EȺ   �    H��I��H��t������H���H�E�H�E�H�E��   �    H��I��H��t������H���H�E��@   H�E��     H�U�H�E�H��H��H�$������H��ЉE��}� t_H�      H�H��I��H�ö������H���H�E�H��I��H�ö������H���H�E�H��I��H�ö������H��и�����-  H�E�H�U�H�M�H�E�H��H��H�v$������H��ЉE��}� u_H�      H�H��I��H�ö������H���H�E�H��I��H�ö������H���H�E�H��I��H�ö������H��и�����  H�EȋU��P,H�EȋPH�Eȋ@ЉE�H�EȋP,H�Eȋ@ �ЋE�ЉE��    I��H�'�������H���H�E�H�E��    �    H��I��H��t������H��ЋU�H�Eȋ@ H�M��	��H�M���H�������H��ЉE��E�    �E�    �   �E���Hc�H�E�H�H�E��E�;�l���}~H�E��@a��ta�E���Hc�H��p���H�H�E���   H��H��I��H�1t������H��ЋE���Hc�H��p���H�H��H��������H��ЃE����E��}�?�e�����H�E�H��I��H�ö������H���H�E�H��I��H�ö������H���H�E�H��I��H�ö������H��ЋE�H�Đ   [A_]���UH��AWSH��`��H�����I���      L�H�}�H�u�H�U�H�M�D�E�H�E�H�E�H�Eغ�   �    H��I��H��t������H���H�E�H��H� ������H���H��H�E�H��H��I��H�:w������H����E�    �"H�U؋E�H����uH�U؋E�H�� �E��}�_~�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉEп    I��H�'�������H���H�E�H�EȺ    �    H��I��H��t������H��ЋU�H�E��@ H�M��	��H�Mȉ�H�������H��ЉEă}� t!H�E�H��I��H�ö������H��ЋE���  �E�    �$�E���Hc�H�E�H�H�E�H�E��@a��t�E��}�?~���H�E��@a���G  �}�?�=  �U�H�E؉PsH�E��@a��E���H�E؈PbH�U�H�E�H��H��H�l!������H���H�U؉BkH�E؋@k���uOH�E�H��H�D�������H�<I�߸    H�r�������H���H�E�H��I��H�ö������H��и   ��   �E���@��t$H�E؋@kH�U�H�M�H�Ή�H�/#������H���H�M�H�E຀   H��H��I��H�1t������H��ЋU�H�E��@ H�M��	��H�Mȉ�H�`������H��ЉEĐH�E�H��I��H�ö������H��и    �JH�E�H��I��H�ö������H���H�E�H��H�h�������H�<I�߸    H�r�������H��Ҹ����H��`[A_]���UH��AWSH��P��H�����I�B�      Lۉ}�H�u�H�U��    I��H�'�������H���H�E��E�    �E��E��E������E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E��E܋E�;E���   �}� tV�E�H�U����H�U�H��H�¾   H�`������H��ЉẼ}� t#H�E�H��I��H�ö������H��и�����?  �E�H�U����H�U�H��H�¾   H�������H��ЉẼ}� t#H�E�H��I��H�ö������H��и������   �E��E�E��E��E�   H�E��@�����E�    ��U�E�EȋE�H��    H�E�HЋ �E�E�H��    H�E�H��     �}��uL�E�H�U����H�U�H��H�¾   H�`������H��ЉE̐H�E�H��I��H�ö������H��ЋE��6�E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��Y���H��P[A_]���UH��AWSH��   ��H�����I���      L�H��h����   I��H�'�������H���H�E�H�E�H�E�H�E�H   H�E�H��h���H�E�H��H��I��H�fS������H���H�U�H�E�H��H��I��H�V������H��п   I��H�'�������H���H�E�H�E��   �    H��I��H��t������H���H��p���H�E�H�E��   �    H��I��H��t������H���H�E��@   H�E��     H�U�H�E�H��H��H�$������H��ЉE�}� t<H�E�H��I��H�ö������H���H�E�H��I��H�ö������H��и    ��  H�E�H�U�H�M�H�E�H��H��H�v$������H��ЉE��}� u<H�E�H��I��H�ö������H���H�E�H��I��H�ö������H��и�����d  H�E��U��P,H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE��    I��H�'�������H���H�E�H�E��    �    H��I��H��t������H��ЋU�H�E��@ H�M��	��H�M���H�������H��ЉE�}� tSH�E�H��I��H�ö������H���H�E�H��I��H�ö������H���H�E�H��I��H�ö������H��ЋE��l  �E�    �   �E������E���Hc�H�E�H�H�E�H�E��@a��t!H�E�H�U�H��H��H�� ������H��ЉE�}� u9H�E��@a �U�H�E��@ H�M��	��H�M���H�`������H��ЉE�}� ��E��}�?�k����}� tPH�E�H��I��H�ö������H���H�E�H��I��H�ö������H���H�E�H��I��H�ö������H��ЋE��uH�E��@kH�U�H�M�H�Ή�H��@������H��ЉE�H�E�H��I��H�ö������H���H�E�H��I��H�ö������H���H�E�H��I��H�ö������H��ЋE�H�Đ   [A_]���UH��H����H�5����I���      Lމ}�E�E��}� u�E��   �E����rH�P     H�H�P     H�����UH��H����H�����I�7�      L�H�}��   H�E�H���r�����UH��AWH����H�����I���      L�H�@     H�H�U�H�H     H�    H�        �    H�M�   �    H��I��H��t������H��ѐH��A_]���UH��AWSH��P��H�����I�t�      Lۉ}��u��}� u
�    ��  H�H     H�H=�   v%H���������H�<I�߸    H�r�������H��ҐH�        ���u�H�        ��PH�        ��E����E�E�%�  ��t�E��E�    �E�    �E�    �}� t�E��   �E�   �K  �}��  �=  H�@     H�H�E�H�E�    �E�    �  H�E؋@����   H�E؋@9E���   H�E�H�H�E؋@��H�H�E�H�E؋@+E���H�E؉PH�E؋P�E��H�E؉PH�E�H�E�H�@     H�H�E��E�    �mH�E؋@��tH�E��E��WH�E�H�E�H�E�H�E�H�E�H�@H�PH�E�H�PH�E��@   H�E�H�U�H�H�E��U��PH�E�H�U�H�P�E���!�}��   ~��H�E��E��}��   ������E�   ���}� ��   H�@     H�H�E��E�    �~H�E؋@��tH�E��E��hH�E�H�E��E��H�\G������H���H�E�H�E�H�U�H��E��E���H�E��PH�E��U��P�E���+E���H�E��PH�E�H�@   ��}��   �u���H�        �    H�H     H�H�PH�H     H�H�E�H��P[A_]���UH��SH��(��H�����I�O�      L�H�}�H�}� ��  �H�        ���u�H�        ��PH�        �H�E�H�E�H�@     H�H�E��E�    �M  H�E�H� H9E�tH�E��E��2  H�E�H�E�H�H     H�H�P�H�H     H�H�E؋@��uH�E�H��H��G������H����   H�E؋@��uH�E�H�@H�E�H�E�H�@H�P�H�E�H�PH�E�H�@H��tH�E؋@����   H�E�H�@H��uRH�E�H� H��H��G������H���H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    ��}��   �������H�        �    ��H��([]���UH��AWH��H��L�����I�M�      M�H�}��u�H�E�    �E�    H�}� u�E��   ��H�}H������I� ���8  �H�        A� ��u�H�        A� �PH�        A� H�@     I� H�E�H�E�H�E��E�    �   H�E�H� H9E�t
H�E��   H�E�H�E��E�   H�E��P�E��=   v@H�H     I� �U�H�E�H��H���������I�< M�Ǹ    I�r�������M�A����H�E�H� H�E�H�E��P�E��H�E��P�E��}��   �X���H�        A�     �}� u�E��   ��H�}H������I� ���H�E�H��HA_]���UH��H�� ��H�����I���      L�H�}�H�u��E�    H�E�H�E��   H�E�� ��H�E��@9�sH�E��P#H�E��@9�rH�E��@#    H�E�f�   H�E�H�PH�E��@#��H�H�E�H�PH�E�H�PH�U�H�U�H�R� �H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  �E��}��E����E�����UH��H�� ��H�����I���      L�H�}�H�u��E�    H�E�H�E�H�E��@'�PH�E��P'H�E��P'H�E��@9�rH�E��@'   �H�E��P#H�E��@'9�r�H�E��@'�P�H�E��P'�JH�E�H�PH�E��@'��H�H�E�H�PH�E�H�PH�E�H�HH�M���H�E��@'�PH�E��P'�E��}�~��E�����UH��AWSH��0��H�����I�Ʈ      L�H�}�H���������H�H� H�E�H�E�H�E�H�E�H��I��H�z������H��ЉE�H�E�H��I��H�z������H��ЉE؋U܋E��=   ~
������   H�E�� </uH�E��E�H�HE�H�m�H�E�� </tH�E�H�E�H�PH�U�� /�H�E�H�U�H�E�H��H��I��H�:w������H���H�E�H��I��H�z������H��Љ�HE�H�m�H�E�� </u	H�E��  �H�E�H�E��  �    H��0[A_]���UH��AWSH����H�����I�w�      L�H���������H�H� H��I��H�z������H��Ѓ�w
�    �   H���������H�H� H�E�H�E�H��I��H�z������H��Љ�HE��H�E�H�P�H�U��  H�E�� </u�H���������H�H� H��I��H�z������H��Ѓ�vH�E��  �    H��[A_]���UH��AWSH��0��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
�    ��  H�E�H��I��H�z������H��ЉE�E�H�H�P�H�E�H�� </u�E�H�H�P�H�E�H��  �}� 
�    �  �}���   H�E�H��� <:u%H�U�H�E�H��H��I��H�:w������H����K  H�$�������H�<I��H���������H���H��H�E�H��H��I��H�:w������H���H�E�H��I��H�z������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H�:w������H����   H�$�������H�<I��H���������H���H��H�E�H��H��I��H�:w������H���H�E�H��I��H�z������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H�:w������H���H�E�H��0[A_]���UH��H����H�����I�K�      L�H�}�H�E�H�E�H�}� u�    �+�E�    �H�E�� </u�E�H�E�H�E�� ��u�E�����UH��AWSH��0��H�����I�ݩ      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
������   H�E�H��I��H�z������H��ЉE�E�H�HE�H�m��H�E�� </tH�m�H�E�� ��t�E�P��U�����H�E�H�U�H�E�H��H��I��H�:w������H���H�E��  �    H��0[A_]���UH��H��0��H�����I���      L�H�}�H�u��U܉M�L�E�H���������H�H� H�E��E�H9E�}?H�E��@��H9E�}0H�E�H�E��E�H�E�H��H�E�H�H��    H�E�HE؉������UH��SH��@��H�����I�a�      Lۉ}ԉuЉỦM�L�E�L�M�f�E�  H�E�H�@H�E�H�E��@�E�}�u�E�    �E�    �   f�E� H�E��@�EȉE��H�H� H�E�H�� f�E�H�E�� ���E��J�E�f#E�f��t5�UЋE��Hc��UԋE��H�H�}��M�U�I��H��H��V������H���f�e�m��}� y��E�H�E��@9E��b�����H��@[]���UH��AWSH��0��H�����I�J�      Lۉ}܉u؉UԉM�D�E�L�M��E�    �X�E�    �CH�E�L��   �M�H�E��P�u؋E��Hc��}܋E��H�H��I��H��V������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I���      Lۉ}܉u؉UԉM�D�E�L�M��E�    �p�E�    �[H�E�H��   �E��E�i��E��A��H�E��P�M؋E��Hc��M܋E��H�I��D��H��I��H��V������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I�ԥ      Lۉ}܉u؉UԉM�D�E�L�M��}� �[  �}� �Q  �E�    �>H�E�L��   �M�H�E��P�E�Hc��}܋E��H�H��I��H��V������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E����Hc��}܋E��H�H��I��H��V������H��ЃE��E�;E�|��E�    �AH�E�H��   �M�H�E��P�u؋E��Hc��E�H�I��H��I��H��V������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E��Hc��}܋E����H�H��I��H��V������H��ЃE��E�;E�|���H��0[A_]���UH��AWSH��@��H�����I�*�      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}��  �E�    ��   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��   �E�f#E�f��tDH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H��V������H����BH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H��V������H���f�e�m��}� �[����E�H�E��@9E��	�����H��@[A_]���UH��SH��8��H�����I�¢      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H��[������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I��      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}���   �E�    �   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��W�E�f#E�f��tBH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H��V������H���f�e�m��}� y��E�H�E��@9E��T�����H��@[A_]���UH��SH��8��H�����I��      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H��]������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I�)�      L�H�}ȉuĉU��M�D�E�D�M�H���������H�H� H�E�H�E�H   � �? �    H��I��H��t������H����E�    �U�H�E��P4�UH�E��P8�UH�E��P<H�E��@H   H�E��@L   H�E��P<H�E��PP�UH�E��PTH���������H�H��H�E�H�PXH�E��@D    H�E��PDH�E��P@�U�H�E��P�U�H�E��P�U�H�E��P �U�H�E��P�U H�E��P`�} u�E�   H�E��@�P�H�E��P(H�E��P�E�)ЍP�H�E��P$H�E��@0   �E����H�E��P,H�E��@��H�E��@��H�E�I���Ѻ    �    I��H�ip������H���H�E��@4��H�E��@����H�E�I��A�ȹ   �   �   H��X������H��Ѓ}� u:H�E��@����H�E�I��A���� �   �   �   H��X������H����8H�E��@����H�E�I��A���� �   �   �   H��X������H��Ѓ}� t}H�E��@����H�U��E�I��A���� ����   �   H��X������H���H�E��@4��H�E��@���ƋE��H�U�I��A�ȹ   ��ƿ   H��X������H���H�E��@8A��H�E��@$��H�E��@(��H�E��@,��H�E��@0��H�E�I��H��X������H���H�E�H��I��H�z������H������E�H�E�H�pHH�E��@��E܉������)Љ�H�E�H���u�I��A���� ������   ��H��H�_������H���H��H�E��@����H�E�I��A�    �   �   �   H�Z������H���H�E�H�PHH�E��@��H���u�I��A���� ������   �ƿX   H��]������H���H��H�E�H�PHH�E��@��(H���u�I��A���� ������   �ƿ-   H��]������H���H��H�E�H�e�[A_]���UH��AWSH��0��H�����I���      L�H�}�H�u�H�E��P0H�E��@Ѓ�P�E�H�E��P,H�E��@Ѓ��E��E�P   �E�   �E�    �E���� H�E�H��I��H�z������H��ЉE�H�E�L�@H�M؋U܋E���������p��E�<�E��������ƋE���)ƋE��H�E�H���u�M��A�ȉщ�H��H�1]������H���H���H�e�[A_]���UH��H����H�����I���      L�H�}��   H�E�H���r�����UH��H����H�����I�h�      L�H�}������UH��H����H�����I�=�      L�H�}�H�U��BD    H�U��JDH�U��J@H�U��R8A��H�U��R$��H�U��R(A��H�U��R,��H�U��R0��H�U�I��D��I��X������J��А����UH��SH��(��L�����I���      Mډ�f�E�H���������I�H� H�E�H���������I�H��H�E�H�PXH�E�@(�P�H�E�@H���к    ��E�H�E�@$�P�H�E�@L���к    ��E�H�E�P<H�E�PPH�E�PD�E�9�rH�E��@D    H�E�@@�PH�E�P@H�E�P@�E�9�r9H�E��@D    H�E�PDH�E�P@H�E�H��H��e������I����E��  f�}���   H�E�@D����   H�E�@D�P�H�E�PDH�E�H�xHH�E�pTH�E�@PH�U�J,H�U�RLA��H�U�R@A��ʃ���H�U�J0H�U�RHA��H�U�RDA��ʃ�A��H���u�I��A������D�޿    H��[������I���H����   f�}�	uH�E�@D�PH�E�PD��   f�}�
u!H�E��@D    H�E�@@�PH�E�P@�   f�}���   H�E�H�xHH�E�pTH�E�PPH�E�H,H�E�@LA��H�E�@@A��ȃ���H�E�H0H�E�@HA��H�E�@DA��ȃ�A���E�H���u�I��A���щ�D�މ�H��[������I���H��H�E�@D�PH�E�PD�E�H�]�����UH��H����H�����I��      L؉}�H���������H�H� H�E��U�H�E��P<�����UH��SH��(��H�����I���      L�H�}�H�}� t=H�E�H�E��&H�E�H�PH�U�� f�����H�Df������H���H�E�� ��u���H��([]���UH��AWSH��P��H�����I�)�      L�H�}��u��U��M�L�E�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H�(�������H�<I�߸    H�r�������H��Ҹ�����6  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H�6�������H�<I�߸    H�r�������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�N�������H�<I�߸    H�r�������H��Ҹ   ��   �E�    �   �E�    �   �}� tNH�E�H��   H�E��P�M��E���E��Hc��M��E���E��H��M�I��H��I��H��V������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H��V������H��ЃE��}� �U����E��}� �;����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��P��H�����I�G�      L�H�}��u��U��M�D�E�L�M�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H�(�������H�<I�߸    H�r�������H��Ҹ�����3  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H�6�������H�<I�߸    H�r�������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�N�������H�<I�߸    H�r�������H��Ҹ   ��   �E�    �   �E�    �   �}� tKH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H��V������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H��V������H��ЃE��}� �X����E��}� �>����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��0��H�����I�d�      Lۉ}܉u؉U�H�M��E�    �   �E�    �t�U�������E��H���������H�Hڋ��E�}� tBH�E�H��   H�EȋP�MԋE��Hc��M؋E��H��M�I��H��I��H��V������H��ЃE��}�~��E��}��o�����H��0[A_]���UH��AWSH��@��H�����I���      Lۉ}̉uȉUĉM�L�E��E���� �E�``` �E���� �EĉE��ẺE܋E��E؋EȉEԋE؍P��E��xH�M��E�I��A�    �   ��I��H�Z������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H�Z������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H�Z������H��ЋEԍP��E܍pH�M��E�I��A�    �Ѻ   ��I��H�Z������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H�Z������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H�Z������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H�Z������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H�Z������H��ЋEԍP��E܍p�M��E�ȃ�H�M�I��A�    �Ѻ   ��I��H�Z������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H�Z������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H�Z������H��ЋE؍P��M܋E�ȍp��E���H�M�I��A�    �   ��I��H�Z������H��АH��@[A_]���UH��H��8��H�����I�Y�      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �CH�E�H�PH�U�� ���E�H�E�H�PH�U�� ���E�E�+E�E�}� u�}� t
�m��}� u��E�����UH��H��8��H�����I�Ë      L�H�}�H�uЉŰẺE�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M����E��P��U���u�H�E�����UH��H�� ��H�����I�L�      L�H�}���U��E�E��E�H�E�H�E��H�E�H�PH�U��U��m��}� u�H�E�����UH��AWSH��0��H�����I��      L�H�}�H�u�H�E�H�E�H�E�H�E��E�    H�E�H�PH�U�� ����I��H�J�������H��ЉE�H�E�H�PH�U�� ����I��H�J�������H��ЉEԋE�+EԉE܃}� u�}� t뗋E�H��0[A_]���UH��AWSH����H�����I�,�      L�H�}�H�u�H�E�H��I��H�z������H��Љ�H�E�H�H�E�H��H��I��H�:w������H���H�E�H��[A_]���UH��H�� ��H�����I���      L�H�}�u�H�E�H�E��H�E�� ��9E�uH�E��H�E�H�E�� ��u۸    ����UH��H�� ��H�����I�T�      L�H�}�H�u�H�E�H�E�H�E�H�E��3H�E��H�E�� 8�u!H�E�� ��H�E�� ��Ѕ�u�    �'H�E�H�PH�U��H�E�H�PH�U�� 8�t����������UH��H��0��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E��  H�E�����UH��AWH��(��H�����I�=�      L�H�}؉uԋU��҉Uԃ}� uOH�U�H��I��H�z������H��҉�H�E�H���   H�E�� ��tH�E�� ��9E�u	H�E��   H�E�H�E؃�H��űE�i��E�H�E�H�E��H�E�H�E� ������H�E� ��!�%������u%H�E� 3E䍐����H�E� 3E���!�%������t�H�E�H�E��H�E�H�E�� ��tH�E�� ��9E�u�H�E�H��(A_]���UH��H��@��H�����I��      L�H�}�H�u�H�U�H�U�H�U������   H�U�H�������   H�E�    H�E�    H�E�    H�E�    �H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�t�H�E�H+E��'H�U����H�Uȉ�H��H��w������H���H+E�����UH��H����H�����I�ޅ      L�H�}�H�E�H�E��H�E�H�E�� ��u�H�E�H+E�����UH��AWSH��@��H�����I���      L�H�}�H�u��U�H�E�H�E�H�E�H�E��E�    �kH�E�H�PH�U�� ����I��H�J�������H��ЉE�H�E�H�PH�U�� ����I��H�J�������H��ЉEԋE�+EԉE܃}� u�}� t
�m��}� u��E�H��@[A_]���UH��H��(��H�����I�ʄ      L�H�}�H�u��U�H�E�H�E�H�E�H�E��}� u)������2H�E�H�PH�U��H�E�H�PH�U�� 8�u�m��}� u����E�����UH��H��8��H�����I�J�      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �!H�U�H�BH�E�H�E�H�HH�M����E��E�9E�w�H�E��  �E�����UH��AWH����H�����I�˃      L�H�}�H�u�H�M�H�U�H��H��I��H��x������H��҉�HE�H�E�� ��tH�E���    H��A_]���UH��AWH��(��H�����I�Y�      L�H�}؉u�H�U�H��I��H�z������H��҉E��U�H�E�H�H�E��E�    �H�E�� ��9E�uH�E��H�m��E��E�9E�wڸ    H��(A_]���UH��H��0��H�����I�Ȃ      L�H�}�H�u�H�E�H� H�E�H�}� u�    �vH�E�H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u,�}� u
H�E�    �H�E�H���  H�E�H�U�H�H�E���}� u������UH��H��@��H�����I��      L�H�}�H�u�H�E�H�E�H�E�    H�E�    H�E�    H�E�    H�E�� ��u
�    ��   H�E�H��� ��u+�H�E�H�E��H�E�� 8�t�H�E�H+E��   H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�u�H�E�H+E�����UH��H��8��H�����I�؀      L�H�}�H�u�H�U�H�}� uH�E�H� H�E�H�}� u
�    ��   �H�E�H�PH�U�� ���E�H�E�H�E��
�E�;E�u��H�E�H�PH�U�� ���E��}� uۃ}� uH�E�H�     �    �   H�E�H��H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u4�}� u
H�E�    �H�E�H��H�E�H�E��  H�E�H�U�H�H�E���}� u������UH��H����H�����I��      L�H�}�H�u�H�u�H�M�H�(       H�H��H�������H�������UH��AWSH�� ��H�����I�G      L�H�}�H�u�H�E�H��I��H�z������H��ЉE��2�U�H�M�H�E�H��H��I��H��s������H��Ѕ�uH�E��H�E�H�E�� ��uø    H�� [A_]���UH��AWSH�� ��H�����I��~      L�H�}�H�E�H��I��H�z������H��Ѓ��E�E��I��H�'�������H���H�E�H�}� u�    �$�U�H�M�H�E�H��H��I��H�1t������H��АH�� [A_]���UH��H��8��H�����I�~      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��U�H�E�H�H�E�H�E�H;E�v[H�E�H;E�sQH�E�H�E��E�HE��H�m�H�m�H�E��H�E��H�E�H;E�u��'H�U�H�BH�E�H�E�H�HH�M���H�E�H;E�u�H�E�����UH��AWH����H�����I�N}      L�H�}�H�u�H�M�H�U�H��H��I��H��v������H���H��A_]���UH��AWH����H�����I��|      Lډ}�H�h�������H�<I�׸    H�r�������H�������UH��H����H�����I��|      L؉}��U���H���������H�Hc��������t�E� �E�����UH��H����H�����I�U|      L؉}��U���H���������H�Hc��������t�m� �E�����UH��AWSH��0��H�����I��{      L�H�}ȉuĉU��M��U�H�E�H��H���������H�<I�߸    I�r�������I�A��H�E�H��I��H���������H���H�E�H�E� �E�H�E� 9E�u��H��0[A_]���UH��AWSH�� ��H�����I�[{      L�H�}�H�u�H�E�� ��u�    �LH�E�� <wuH�E�H��I��H��������H���H�U�H�E�H��H��I��H�Z������H���H�E�H�E�H�� [A_]���UH��AWH����H�����I��z      L�H�}�H�U�H��I��H��������H���H��A_]���UH��AWH����H�����I�{z      L�H�}�H�U�H��I��H��������H���H��A_]���UH��AWH����H�����I�0z      L؉}�H�u�H�M��U�H�Ή�I��H�#������H���H��A_]���UH��AWSH�� ��H�����I��y      L�H�}�H�}� u������VH�E�H��I��H�?������H��ЉE�H�E؋@��u+H���������H�H��E�H�։�I��H�#������H��ЋE�H�� [A_]���UH��AWH����H�����I�Ey      L؉}�H�u�H�M��U�H�Ή�I��H�������H���H��A_]���UH��AWH����H�����I��x      L�H�}�H�U�H��I��H��������H���H��A_]���UH��AWSH��@��H�����I��x      L�H�}ȉu�H�U�H�}� u	H�E��  H�E�H�E�H�E�H�E��E�    H�E�H��I��H�?������H��ЉEԃ}����   H�E��@��u7�}�u�}� ~+H���������H�H��E�H�։�I��H�#������H��Ѓ}�
tk�E�;E�}E�}�u�}� ~H�E�H;E�vH�m��m��:�}��^���H�E�H�PH�U�UԈ�E��D����}�u�}� ~�m���E��)�������}�~	H�E��  ��Eԉ�H�E�H�E�H��@[A_]���UH��AWSH�� ��H�����I�Kw      L�H�}�H�u�H�}� u�    �^�E�    �2�E�Hc�H�E�H�� ��H�U�H�։�I��H�������H��ЃE�H�E�H��I��H�z������H��ЋU�9�w��E�H�� [A_]���UH��AWH��(��H�����I��v      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I�������I�A��H��(A_]���UH��AWH��(��H�����I�Kv      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I��������I�A��H��(A_]���UH��AWH����H�����I��u      L�H�}�H�U�H��I��H��B������H���H��A_]���UH��AWH����H�����I��u      L�H�}�H�U�H��I��H��������H��ҐH��A_]���UH��AWH��(��H�����I�Wu      L�H�}�H�u��U܋U�H�u�H�M�H��I��H��������H���H��(A_]���UH��H����H�����I� u      L�H�}�H�}� u������!H�E��P#H�E���+  9�r�������    ����UH��AWH����H�����I��t      L�H�}�H�U�H��I��H�a������H���H��A_]���UH��AWSH��`  ��H�����I�Vt      L�H������H������H�������E�    �E�    �  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H�)�������H���	E�}���  �E�H��    H�h  H�H�h  H�>��H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E��E�H������H�։�I��H���������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�}� t(H������H�E�H��H��I��H���������H����O  H������H��H���������H�<I��H���������H����   H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E�H�������E�H�։�I��H�k�������H���H������H������H��H��I��H���������H����w  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������
   H��H��I��H���������H���H������H������H��H��I��H���������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������   H��H��I��H���������H���H������H������H��H��I��H���������H����  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�EȾ   H��fHn�I��H���������H���H������H������H��H��I��H���������H����]  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eк
   H��H��I��H�=�������H���H������H������H��H��I��H���������H����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ
   H��H��I��H���������H���H������H������H��H��I��H���������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ   H��H��I��H���������H���H������H������H��H��I��H���������H����G  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�E�   H��fHn�I��H���������H���H������H������H��H��I��H���������H����   H������H�ƿ%   I��H���������H��ЋE�Hc�H������H�� ��H������H�։�I��H���������H����4�E�Hc�H������H�� ��H������H�։�I��H���������H��ЃE��E�Hc�H������H�� ��������    H��`  [A_]���UH��H����H�����I��k      L؉��E��E�    �E��S��%wa��H��    H��`  H�H��`  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I�k      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��H�� ��H�����I�6j      L�H�}�H�u�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E�����UH��AWSH��  ��H�����I��i      L�H������H������H��x����E�    H������H�E�f�E�  �E� �E�    �/  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H���������H���	E܃}���  �E�H��    H�r_  H�H�g_  H�>��H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E��E�H�U�H�E�H��H��H���������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H�}� t'H�U�H�E�H��H��H���������H���H�E��e  H�E�H���������H�4H��H���������H���H�E��7  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E�H�������E�H�։�I��H�k�������H���H������H�E�H��H��H���������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������
   H��H��I��H���������H���H������H�E�H��H��H���������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������   H��H��I��H���������H���H������H�E�H��H��H���������H���H�E��3  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�E��   H��fHn�I��H���������H���H������H�E�H��H��H���������H���H�E��x  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�E��
   H��H��I��H�=�������H���H������H�E�H��H��H���������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ
   H��H��I��H���������H���H������H�E�H��H��H���������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ   H��H��I��H���������H���H������H�E�H��H��H���������H���H�E��e  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�Eо   H��fHn�I��H���������H���H������H�E�H��H��H���������H���H�E��   H�E�H���������H�4H��H���������H���H�E�fǅ����  �E�Hc�H������H�� ������H������H�E�H��H��H���������H���H�E��8�E�Hc�H������H�� �E�H�U�H�E�H��H��H���������H���H�E��E��E�Hc�H������H�� �������H�E��  H�U�H������H)�H��H�Ā  [A_]���UH��H����H�����I��`      L؉��E��E�    �E��S��%wa��H��    H�X  H�H�	X  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I�F`      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H�*�������L��Љ�<�����<���Hc�H�����H��  ��<���H���   A_]���UH��AWH���   ��L�����I�E_      M�H����������H�����H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H����������H�����H��M��H���������L��Љ�<�����<���H���   A_]���UH��AWSH��0��H�����I�Z^      L�H�}؉u�H�U�H�M��}�   v
�    �   H�U�H�E�H��H�@       H�<I��H�*�������H��ЉE�}���  ~�   �I�E�E�}� ~:�U�H�E�H�@       H�4H��I��H�1t������H��ЋE�Hc�H�E�H��  �E�H��0[A_]���UH��AWH����H�����I��]      L؉}�H���������H�H�
�U�H�Ή�I��H�������H���H��A_]���UH��AWSH�� ��H�����I�%]      L�H�}�H�}� tj�E�    �?H���������H�H��E�Hc�H�E�H�� ��H�։�I��H�������H��ЃE�H�E�H��I��H�z������H��ЋU�9�w���H�� [A_]���UH��AWH���   ��L�����I�}\      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I��[      M�H��8���H��0���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�H���������I�<M�׸    H�r�������L�������UH��AWH����H�����I��Z      L�H�}�H�U�H��I��H�̢������H��ҐH��A_]���UH��AWH��(��H�����I��Z      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H�K�������H��Ѹ    H��(A_]���UH��AWH��(��H�����I�9Z      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H�K�������H����H�E�H�E�� < tH�E�H   H9E�sH�E�� <
u�H�E��  H�E�H;E�����H��(A_]���UH��AWSH��0��H�����I��Y      L�H�}�H�uЉỦM�H�@      H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H�K�������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H�@      H�H�E�H�@      �0H�@      �D �}�u-�U�H�E�    H��I��H��������H���H�U�H��   �}�u+�U�H�E�    H��I��H�>�������H��Љ�H�EЉ�[�}�u,�U�H�E�    H��I��H�>�������H��Љ�H�E�f��)�U�H�E�    H��I��H�>�������H��Љ�H�EЈ�    H��0[A_]���UH��AWSH��0��H�����I��W      L�H�}�H�uЉỦM�H�@     H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H�K�������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H�@     H�H�E�H�@     �0H�@     �D �}�u'H�E�H��I��H���������H����Z�H�E�� �+�}�u%H�E�H��I��H���������H���fH~�H�U�H��    H��0[A_]���UH��SH��8��H�����I��V      L�H�}�H�u�H�U��E�    �E�    ��  �E�    �E�Hc�H�E�H�� ������%��  �E��E�Hc�H�E�H�� ������lu�E��E�   �E�Hc�H�E�H�� ����H���������H���	E�}��o  �E�H��    H��N  H�H��N  H�>��H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H�T�������H�����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H���������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�[�������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�[�������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H����?  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�[�������H�����   H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�[�������H����jH�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H������E��E�Hc�H�E�H�� ��������E�H��8[]���UH��H����H�����I�\R      L؉��E��E�    �E��S��%wa��H��    H��K  H�H�xK  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��Q      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H�<�������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I��P      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H�<�������L��Љ�<�����<���H���   A_]���UH��H����H�����I��O      L؉}�H�u�H�}� u������w�}��u������jH�E��@#��tH�E��@#�P�H�E��P#H�E��@#H�U��J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U���E�����UH��AWSH����H�����I�O      L�H���������H�H� H��I��H�?������H��ЉE�}��t+H���������H�H��E�H�։�I��H�#������H��ЋE�H��[A_]���UH��AWH��(��H�����I��N      L�H�}�H�u�H�U�H���������H�<I�ϸ    H�r�������H�������UH��H����H�����I�:N      L�H�}��	   H�E�H���r�����UH��SH����H�����I� N      L�H�}�H�}� u.H�@     H�<H���������H���H�@     H��H�E�H��H���������H���H�E�H��[]���UH��AWSH��0��H�����I�~M      L�H�}�H�u�H�E�H���������H�4H��I��H���������H���H�E�H�}� u
������   �E�    H�E�H��I��H�z������H��ЉE܃}�`~	�E�   �$H�E�H�P+H�E�H��H��I��H�:w������H���H�E��@���H�E��PH�E�H��I��H�,�������H��ЋE�H��0[A_]���UH��H��0��H�����I��L      L؉}�H�u�H�E�H�E��E܉E��E�    �}� y,H�E�H�PH�U�� -�}�   �u�E�����E���E��؉E�H�E�H�E�M�Hc�Hi�gfffH�� ��������)�����)��ʉЍH0H�E�H�PH�U�ʈ�E�Hc�Hi�gfffH�� ����)ЉE�}� u��}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWSH��@��H�����I�?K      L�H�}�H�u��U�H�}� u#H�E�H�E�H�E�H�PH�U�� 0H�E��  �  H�E�H�E؋E�Hc�H�E�H�H�E��3H�E؃��E�H�m��}�	~�7   ��0   �U��H�m���H�E�H�E�H;E�wËE�Hc�H�E�H��  H�E�H�E��E�    �8H�E�� <0uH�E��"H�U�H�E�H��H��I��H�:w������H�����E��E�;E�|�H�E�H�E�H�E�H��I��H�z������H��Љ�H�E؋E�H�U�)Љ�H�M�H�E�HȾ    H��I��H��t������H���H��@[A_]���UH��AWH����H�����I��I      L؉}�U�    ��I��H�}H������H���H��A_]���UH��AWH����H�����I�~I      L؉}�u�U��U��I��H�'�������H���H��A_]���UH��AWH����H�����I�/I      L�H�}�H�U�H��I��H��K������H��ҐH��A_]���UH��AWH����H�����I��H      L�H�}�u�M�H�U��H��I��H��M������H���H��A_]���UH��H����H�����I��H      L؉}�u�E��}�E��E��}�ЉE��}� x�E���y�E����E��E�+E�E��!�}� y�E���~�E����E��U��E�ЉE�H�E�����UH��H�� ��H�����I�
H      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H�� ��H�����I�`G      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H��H��H�����I��F      L�H�}�H�u��U�H�E�H�E�H�E�H�PH�U�� ���E�E���H���������H�H������ ��uǃ}�-u�E�   H�E�H�PH�U�� ���E��"�E�    �}�+uH�E�H�PH�U�� ���E�}� t�}�u9�}�0u3H�E�� <xtH�E�� <XuH�E�H��� ���E�H�E��E�   �}� u�}�0u�   ��
   �E��}� t	H��   ������H�E�E�Hc�H�E�H�H��H�ЉE؋E�Hc�H�E�H�H��H�E�}� t�}� ~�E�)E�H�E��]�H�E�    �E�    �E���H���������H�H��������t�m�0�[�E���H���������H�H���������5  �E���H���������H�H��������t�7   ��W   )E�E�;E���   �}� ��   �}� tgH�E�H;E�|H�E�H;E�u0�E�;E�~(�E�����H�E�   �H���������H�� �����   �E�   �E�H�H�U�H��H�E��E�H�H)E��eH�E�H;E�H�E�H;E�u-�E�;E�~%�E�����H�E����H���������H�� �����$�E�   �E�H�H�U�H��H�E��E�H�HE���H�E�H�PH�U�� ���E��y������H�}� t�}� t
H�E�H���H�E�H�U�H�H�E�����UH��AWH����H�����I��C      L�H�}�H�M�
   �    H��I��H�>�������H���H��A_]���UH��AWH����H�����I�-C      L�H�}�H�M�
   �    H��I��H�>�������H���H��A_]���UH��AWAVAUATSH����H�����I��B      L�H�}�H�uȉU�L�eп    L��L�`� �؉���H���������H�H������ ��uЃ�-u�   L��L�`� �����+uL��L�`� �؃}� t�}�u-��0u(A�$<xt	A�$<XuI�D$� ��I���E�   �}� u��0u�   ��
   �EċE�Hc������    H��I�ǋE�Hc������    H��H�Љ�A�    A�    ����H���������H�H��������t��0�T����H���������H�H��������tz����H���������H�H��������t�7   ��W   )�;]�}GE��x
M9�wM9�u��9�~A������A�   �E�H�L��Hc�I�L��L�`� ���;������E��yA�����H���������H�� "   �	����tI��H�}� tE��tI�D$��H�E�H�U�H�L��H��[A\A]A^A_]���UH��H����H�����I��@      L؉}��   �   ���r����UH��AWSH����H�����I�T@      L�H�}�H�E�H���������H�4H��I��H��v������H��Ѕ�uH���������H�H� ��    H��[A_]���UH��AUATSH�� ��H�����I��?      L�H�}�H�u�H��     ��E�L�e�H�]�E�,$L��L�`��H��H�XD�(�m��}� uې�H�� [A\A]]���UH��H��8��H�����I�e?      L�H�}�H�u�H�U�H��     ��E�H�E�H�E�H�E�H�E�H�E�H�E�H�E�� ���E�H�E�H�PH�U�H�U���H�E�H�PH�U�H�U���H�E�H�PH�U��U���m��}� u�������UH��SH��H��H�����I��>      L�H�}�H�u�H��     ��E�H�E�H+E��EȋE�9E���  �E�����EȺ    ��E��EȋU�H�E�H�H�E�H�E�H�E�H�E�H�E�E�H�H��H��H�E�H�H�E�H�E�H;E�sjH��     H�H�U�H�E�H��H���щEă}� u/�E�H�H��HE�H�U�H�E�H��H��H��������H�����  �}� y�E�H�HE���  �H�E�H;E���   H��     H�H�U�H�E�H��H���щEă}� u)�E�H�HE�H�U�H�E�H��H��H��������H���뢃}� ��   H�E�H;E�uA�E�H�HE�H�U�H�M�H�E�H��H��H���������H��ЋE�H�HE�H�E�H�E��M���H�U�H�E�H��H��H��������H��ЋE�H�H��HE��E�H�HE���   �E�H�H��HE�����H�E�H;E���   H�E�H+E�H��H�E�H+E�H9�|4�E�Hc�H�E�H�H�E�H��H��H�=�������H���H�E�H�E������H�U�H�E�H��H��H�=�������H��ЋE�Hc�H�E�H�H�E������E�H�H��HE�H�U�H�M�H�E�H��H��H���������H��ЋE�H�H��HE�H�E�H�E������H��H[]���UH��H�� ��H�����I��;      L�H�}��u�U�H�M�H��     H�U�H��U�H��     ��U��U���H�U�H�H�U�H��H��H�=�������H��А����UH��AWH����H�����I�B;      L�H�}�H���������H�<I�׸    H�r�������H��Ѹ����H��A_]���UH��H��@��H�����I��:      L�H�}�H�u�H�U�H�U��H�E�H�U����H���������H�Hc���҃� ��u��E�    H�U���҃�+t��-u�E�   H�E�H�����������E��E�    �E�    �E�    �;�M�H�����������Y�H�U���҃�0�*��X��E�H�E��E�H�U����H���������H�Hc���҃���u�H�U����.uuH�E��?�M�H�����������Y�H�U���҃�0�*��X��E�H�E��E��E�H�U����H���������H�Hc���҃���u��U�)U�}� uH���������f���  �}� t�E�H���������f(fW��E�H�U����etH�U����E��   �E�    H�E�H�U���҃�+t��-u�E�   H�E��E�    �%�M܉����҉�H�U���҃�0ʉU�H�E�H�U����H���������H�Hc���҃���u��}� t�U�)U���U�U�}����|	�}�   ~H� ���������   H�����������E��E�E܃}� yF�]��A�E܃���t&�}� y�E��^E��E���E��YE��E��}��E��Y��E��}� u�H�}� tH�E�H�U�H��E�����UH��H����H�����I��7      L؉}�H�E�   �E�    �H�U�H��H��H�H�H�E��E��E�;E�|�H�E�����UH��AWSH��@��H�����I�Q7      L��E�H�}��u�H�}� u	H�E��  H�E�H�E�H���������f��f/E�v,H�E�H�PH�U�� -�E�H� �������f(fW��E��E�H��������f/s�E��H,�H�E��/�E�H����������\��H,�H�E�H�       �H1E�H�E�H�E�H�E�H��x�H*��H��H���H	��H*��X��M��\�f(��EȋE���H�A�������H���H��x�H*��H��H���H	��H*��X��YE�H��������f/s�H,�H�E��*H����������\��H,�H�E�H�       �H1E�H�E�H�E�H�M�H�U�H�E�H���������H�43H��I�߸    I���������I�A��H�E�H��@[A_]���UH��AWH����H�����I�g5      L�H�}�H�U�    H��I��H��������H���H��A_]���UH��AWH����H�����I�5      L�H�}�H�u�H�M�H�U�H��H��I��H��������H����Z�H��A_]���UH��AWH��(��H�����I��4      L�H�}�H�u�H�M�H�U�H��H��I��H��������H����E��E�H��(A_]���UH��H����H�����I�a4      L؉}��E����3E�)�����UH��H��@��H�����I�-4      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�    H�}� y>H�E�H�PH�U�� -H�       �H9E�uH��������H�E�H�E��H�E�H��H�E�H�E�H�E�H�M�H�gfffffffH��H��H��H��H��?H)�H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U��ʈH�M�H�gfffffffH��H��H��H��H��?H)�H��H�E�H�}� u�H�}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U߈H�E�H;E�w�H�E�����UH��AWH��8��H�����I��2      L�H�}�H�uЉU�H�U�H�U�H�}� yH�U�H�JH�M��-H�]�H�U�H�U��}�u$H�M�H�u�   H��I��H���������H����H�M�H�U�H��H��H���������H���H�E�H��8A_]���UH��H��0��H�����I�2      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E�H�M�H���������H��H��H��H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U�ʈH�E�H���������H��H��H��H�E�H�}� u�H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWH��8��H�����I�1      L�H�}�H�uЉU�H�U�H�U�H�U�H�U��}�u$H�u�H�M�   H��I��H���������H����H�M�H�U�H��H��H���������H���H�E�H��8A_]���UH��H����H�����I�z0      L؉}������UH����H�����I�T0      Lظ   ]���UH��H����H�����I�)0      L�H�}��    ����UH��H����H�����I��/      L�H�}�H���������H�H� ����UH��H����H�����I��/      L�H�}�H���������H�H� ����UH��H�� ��H�����I��/      L�H�}��u�H�U�H�M�    ����UH����H�����I�N/      Lظ    ]���UH��H����H�����I�#/      L��E�H��������f������UH��H����H�����I��.      L��E�H��������f������UH��H����H�����I��.      L��E��}�H��������f������UH��H����H�����I�u.      L��E�H�}�H��������f������UH��H����H�����I�8.      L��E��M�H��������f������UH��H��(��H�����I��-      L��E��M��E��U��U��E��E��E������������������������������]��E�����UH��H����H�����I��-      L��E����E����]��E�����UH��H����H�����I�Q-      L��E�H� �������f������UH��H����H�����I�-      L��E�H�(�������f������UH��H����H�����I��,      L��E�H�0�������f������UH��H����H�����I��,      L��E�H�8���������E��E�����UH��H����H�����I�b,      L��E�H�@�������f������UH��H����H�����I�),      L��E�H�H�������f������UH��H����H�����I��+      L��E�H�P�������f������UH��H����H�����I��+      L��E�H�X�������f������UH��AWH����H�����I�|+      L��E��E�H�`�������H�f(�fHn�I��H���������H���H��A_]���UH��H����H�����I�+      L؉}�H�u�    ����UH��AWH����H�����I��*      Lډ}�H�u�H�h�������H�<I�׸    H�r�������H�������UH��AWH��(��H�����I��*      Lى}�H�u�H�U�H�y�������H�<I�ϸ    H�r�������H�������UH��AWSH�� ��H�����I�<*      L�H�}�H���������H�<I�߸    H�r�������H����E�    �.�E�H�H��    H�E�HЋ ��I��H�p�������H��ЃE��}�?~̸����H�� [A_]���UH��AWH����H�����I��)      L�H�}�u�H���������H�<I�׸    H�r�������H�����f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�                                                                         ~ � � � � � � � � ~             ~ � � � � � � � � ~                 l � � � � | 8                   8 | � | 8                   < < � � �   <                < ~ � � ~   <                      < <              � � � � � � � � � � � � � � � �           < f B B f <           � � � � � � � � � � � � � � � �        2 x � � � � x             < f f f f <  ~               ? 3 ? 0 0 0 0 p � �              c  c c c c g � � �               � < � < �             � � � � � � � � � � �               > � >                  < ~    ~ <                f f f f f f f   f f              � � � {                | � ` 8 l � � l 8  � |                       � � � �              < ~    ~ <  ~              < ~                           ~ <                      �                         0 ` � ` 0                         � � � �                       ( l � l (                      8 8 | | � �                   � � | | 8 8                                                 < < <                  f f f $                             l l � l l l � l l           | � � � |   � � |               � �   0 ` � �             8 l l 8 v � � � � v           0 0 0 `                             0 0 0 0 0 0               0         0                   f < � < f                         ~                                    0                     �                                                           0 ` � �             8 l � � � � � � l 8              8 x       ~             | �    0 ` � � �             | �   <    � |               < l � �                 � � � � �    � |             8 ` � � � � � � � |             � �     0 0 0 0             | � � � | � � � � |             | � � � ~     x                                                       0                  0 ` 0                      ~     ~                     ` 0      0 `             | � �                       | � � � � � � � |              8 l � � � � � � �             � f f f | f f f f �             < f � � � � � � f <             � l f f f f f f l �             � f b h x h ` b f �             � f b h x h ` ` ` �             < f � � � � � � f :             � � � � � � � � � �             <         <                   � � � x             � f f l x x l f f �             � ` ` ` ` ` ` b f �             � � � � � � � � � �             � � � � � � � � � �             | � � � � � � � � |             � f f f | ` ` ` ` �             | � � � � � � � � |           � f f f | l f f f �             | � � ` 8   � � |             ~ ~ Z       <             � � � � � � � � � |             � � � � � � � l 8              � � � � � � � � � l             � � l | 8 8 | l � �             f f f f <     <             � � �   0 ` � � �             < 0 0 0 0 0 0 0 0 <               � � � p 8                 <         <          8 l �                                                   �       0                                     x  | � � � v             � ` ` x l f f f f |                   | � � � � � |                < l � � � � v                   | � � � � � |              6 2 0 x 0 0 0 0 x                   v � � � � � |  � x       � ` ` l v f f f f �                 8      <                        f f <       � ` ` f l x x l f �             8         <                   � � � � � � �                   � f f f f f f                   | � � � � � |                   � f f f f f | ` ` �             v � � � � � |                � v f ` ` ` �                   | � ` 8  � |              0 0 � 0 0 0 0 6                    � � � � � � v                   � � � � � l 8                   � � � � � � l                   � l 8 8 8 l �                   � � � � � � ~   �             � �  0 ` � �                 p                                        p         p                       v �                        8 l � � � �                               ��� ��� ~~~                                 uuu ��� ��� ���                                 ��� ��� ��� ��� ;;;                          ��� ��� ~~~ ��� ���                         ��� ��� ���     ��� ���                         ��� ���      ��� ��� ppp                 @@@ ��� ���         III ��� ���                 ��� ��� ��� ��� ��� ��� ��� ���                 ��� ���                 zzz ��� ���         ``` ��� ���                     ��� ���         ��� ��� MMM                     ��� ��� bbb     ��� ���                         ||| ��� ���      ��C%lf, %lf
             9@      �Entrada maior que o limite
 Erro ao criar o arquivo "%s"
       Error ao criar o arquivo "%s", atingio o limite de arquivos na entrada de directorio
   Panic: __malloc, sem espaco na tabela de alocacao
      panic: realoc sem espaco, %lx size = %d %d
 PWD BitMAP error
 Not suport BitMAP 4-bit Not suport BitMAP > 8-bit strerrorr
              (((((�AAAAAABBBBBB                                �Dubug: %s %x %x
        (null)  Ξ��������������|�������9����������������������@�������@�������Ξ������Ξ������Ξ������Ξ������Ξ������Ξ������Ξ������Ξ������Ξ������Ξ������Ξ����������������������`���������������������0�������f�������f�������f�������f�������K�������f�������f�������f�������f�������f�������f�������f�������f�������f�������f�������'�������9�������f�������]�������T�������f�������9�������f�������f�������f�������f�������f�������f�������f�������f�������f�������0�������f�������B�������f�������f�������K�������(null) %        r���������������*����������������������;���������������������r�������r�������r�������r�������r�������r�������r�������r�������r�������r�������r���������������U�������������������������������������<�������<�������<�������<�������!�������<�������<�������<�������<�������<�������<�������<�������<�������<�������<����������������������<�������3�������*�������<��������������<�������<�������<�������<�������<�������<�������<�������<�������<��������������<��������������<�������<�������!�������panic: sscanf()
        ɴ������}��������������G���������������ɴ��������������������ɴ������ɴ������ɴ������ɴ������ɴ������ɴ������ɴ������ɴ������ɴ������ɴ������ɴ����������������������ɴ������`�������`���������������ʹ������ʹ������ʹ������ʹ��������������ʹ������ʹ������ʹ������ʹ������ʹ������ʹ������ʹ������ʹ������ʹ������ʹ����������������������ʹ������Ĵ��������������ʹ��������������ʹ������ʹ������ʹ������ʹ������ʹ������ʹ������ʹ������ʹ������ʹ��������������ʹ��������������ʹ������ʹ��������������panic: freopen()
 r+ PWD call system funtion error. 
                 $@       �        %lu.%lu                �              �C                                                                        �_�
�@panic: signal()
 panic: sigaction()
 panic: setjmp()  panic: longjmp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �   �  �   �  �   � �    �   � �    �  �   8 �    �  �   � �   H �   h �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          zR x�  ,      @ ���   E�CG����B�A�       $   L   ����    E�CG����B�A�(   t   y��Z   E�CG��G�B�A�      �   ���   E�C�   �   ����    E�C��    �   -���    E�C��        ���p    E�CF�`�A�$   $  ���    E�CG����B�A�$   L  ���r    E�CG��_�B�A�(   t  ��   E�CG��	�B�A�   $   �  ����   E�CF���A�       �  �
���    E�CE���A�    �  ?���    E�CE���A�     ����    E�C��    0  ���A    E�Cx�      P  ���i    E�C`�        t  ���U    E�CL�    �  (��U    E�CL�    �  ]��i    E�C`�    �  ���g    E�C^�    �  ����    E�C�� $     ����   E�CE�{�A�      <  ��9    E�Cp�  $   \  /���    E�CG����B�A�   �  ���^    E�CU� (   �  .��   E�CG���B�A�   (   �  ���   E�CG����B�A�   (   �  ���]   E�CG��J�B�A�   (   (  ���   E�CG��l�B�A�   (   T  9��D   E�CJ��.�B�A�   (   �  Q!��:   E�CG��'�B�A�   $   �  _"��    E�CG����B�A�   �  7#���    E�C��    �  �#���    E�C�� (     �$���   E�CJ����B�A�   (   @  b(��i   E�CG��V�B�A�   (   l  �+��H   E�CG��5�B�A�   (   �  �-��e   E�CJ��O�B�A�      �  �1��a    E�CX�    �  52��9    E�Cp�        N2���    E�CF�w�A�(   (  �2��'   E�CG���B�A�   $   T  �5��   E�CE���A�   $   |  �7���   E�CF���A�      �  �8��    E�C��    �  �9���    E�C�� (   �  �:��O   E�CG��<�B�A�   $     �;���    E�CG����B�A�(   8  �<��C   E�CG��0�B�A�      d  �>��k    E�Cb� $   �  �>���    E�CG����B�A�   �  �?���    E�C�� $   �  "@��   E�CE��A�   $   �  A���    E�CG����B�A�$     �A���    E�CG����B�A�(   D  5B���   E�CG����B�A�   (   p  �C��j   E�CG��W�B�A�       �  �D���    E�CE���� (   �  �E��   E�CG���B�A�       �  |F���    E�CE���� (   	  G���   E�CG��q�B�A�   $   <	  lK��   E�CG����B�A�   d	  KL��9    E�Cp�     �	  dL��+    E�Cb�     �	  oL���    E�C��     �	  �L���   E�CE����   �	  ~O��I    E�C@�     
  �O��u    E�CE�f�A�(   ,
  �O���   E�CG����B�A�   (   X
  �R���   E�CG����B�A�   $   �
  eU���    E�CG����B�A�,   �
  V��2   E�CG���B�A�          �
  Y���    E�C��    �
  �Y��w    E�Cn�      �Y��b    E�CY� $   <  *Z���    E�CG����B�A�$   d  �Z��z    E�CG��g�B�A�   �  [��a    E�CX�    �  P[���    E�C��    �  �[��{    E�Cr� $   �  %\��+   E�CF��A�        (]��6   E�C-�   4  >^��L    E�CC� $   T  j^���    E�CG����B�A�   |  
_���    E�Cw�    �  j_��}    E�Ct� $   �  �_��r    E�CF�b�A�    $   �  `���    E�CF���A�         |`���    E�C��    ,  a��3   E�C*�   L  ,b��7   E�C.�   l  Cc��W    E�CN� $   �  zc���    E�CG����B�A�$   �  �c���    E�CG����B�A�   �  bd���    E�C�� $   �  e��V    E�CF�F�A�       $  2e��P    E�CF�       D  be��U    E�CL�    d  �e��U    E�CL� $   �  �e���    E�CG����B�A�$   �  Ff���    E�CG����B�A�$   �  �f��K    E�CF�{�A�     $   �  �f��K    E�CF�{�A�     $   $  �f��S    E�CF�C�A�    $   L  %g���    E�CG����B�A�$   t  �g��S    E�CF�C�A�    $   �  �g��K    E�CF�{�A�     ,   �  �g��[   E�CG��H�B�A�       $   �  i���    E�CG����B�A�$     �i��]    E�CF�M�A�    $   D  �i��]    E�CF�M�A�    $   l  �i��K    E�CF�{�A�     $   �  j��L    E�CF�|�A�     $   �  ;j��Y    E�CF�I�A�       �  lj��Y    E�CP� $     �j��K    E�CF�{�A�     (   ,  �j���   E�CJ��{�B�A�       X  -s���    E�C��     $   |  �s���    E�CI���A�       �  vt��l    E�Cc� (   �  �t���   E�CJ����B�A�       �  k}���    E�C��     $     �}��   E�CI���A�    $   <  �~���    E�CI���A�    $   d  ����    E�CG����B�A�$   �  @���\    E�CF�L�A�    $   �  t����    E�CG����B�A�$   �  ����    E�CI���A�         �����    E�CI�    $   $  @���L    E�CF�|�A�         L  d���e    E�CF�U�A�    p  �����    E�CF���A�(   �  #����   E�CG����B�A�   (   �  ����=   E�CG��*�B�A�   $   �  ����\   E�CE�M�A�        �����    E�C�� $   4  j����    E�CI���A�    $   \  -����    E�CI���A�       �  �����    E�C�� $   �  �����    E�CG��z�B�A�   �  ���Y    E�CF�       �  *���9    E�Cp�  $     C����    E�CE�q�A�    $   4  �����    E�CG����B�A�   \  k���G   E�C>�,   |  ����u   E�CG��b�B�A�       $   �  א��M    E�CF�}�A�     $   �  ����O    E�CF��A�     $   �  #���L    E�CF�|�A�     $   $  G���S    E�CF�C�A�       L  r����    E�C�    l  ڑ���    E�C��    �  d����    E�C��    �  ���2   E�C)�$   �   ���U    E�CF�E�A�    $   �  -���U    E�CF�E�A�    4     Z���L   E�CM�����-�B�B�B�B�A�      T  n���7    E�C       $   t  ����w    E�CG��d�B�A�(   �  Ԙ��{    E�CI���d�B�B�A�   �  #����    E�C�� $   �  �����   E�CE���A�         {����    E�Cx�     $   4  ؜��\    E�CF�L�A�       \  ���5   E�C,�   |  !���_    E�CV� ,   �  `����   E�CG����B�A�       $   �  ���P    E�CF�@�A�    $   �  C���Z    E�CF�J�A�    $     u���^    E�CF�N�A�       D  ����4    E�Ck�     d  ����v   E�Cm�$   �  ����    E�CF���A�       �  �����    E�C�� $   �  u����    E�CF���A�       �  ���*    E�Ca�       ���'    E�C^�     4  ���/    E�Cf�     T  ���;    E�Cr�     t  ���;    E�Cr�     �  8���:    E�Cq�     �  R���'    E�C^�     �  Y���9    E�Cp�     �  r���9    E�Cp�       ����<    E�Cs�     4  ����=    E�Ct�     T  Ħ��>    E�Cu�     t  ���n    E�Ce�    �  0���;    E�Cr�     �  K���9    E�Cp�     �  d���9    E�Cp�     �  }���9    E�Cp�       ����D    E�C{�     4  ����9    E�Cp�     T  ӧ��9    E�Cp�     t  ���9    E�Cp�     �  ���9    E�Cp�  $   �  ���a    E�CF�Q�A�       �  W���2    E�Ci�     �  i���T    E�CF�     ����X    E�CF�$   4  ݨ���    E�CG����B�A�   \  P���T    E�CF�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            GCC: (Ubuntu 9.3.0-17ubuntu1~20.04) 9.3.0                                        �                  �  �                   �                 ` �                 � �                    �                                     ��                     ��_ cole _             ��                )        �           =         �           0    ��                7    ��                >      x �           C      � �           H      h �           M    ��                T    ��                >      � �           C      � �           H      � �           �   ��                Z     � �          >        �           C      X �           j    ��                q    ��                >      � �           x    ��                ~    ��                �    ��                �    ��                >      � �           C      � �           H      � �           �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                   ��                   ��                   ��                (   ��                2   ��                <   ��                F   ��                O   ��                X   ��                a    � �          k   ��                t   ��                }   ��                �   ��                �   ��                >      � �           �   ��                �   ��                �   ��                �   ��                >      � �           �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                   ��                   ��                   ��                   ��                %   ��                ,   ��                4   ��                ?    ��  �   �       >      � �           5   ��                B   ��                ?    _�  �   �       >      � �           C      � �           C   ��                N   ��                M   ��                Y    � �          `   ��                �   ��                6   ��                j   ��                >      � �           s   ��                |   ��                �    ��  �   e       U    �  �   �       �    ��  �   �      �    � �          �    _�  �   =      �    � �          ?    ��  �   �       }   ��                ~   ��                �   ��                �   ��                �   ��                >      �
 �           �   ��                �    � �   `       �   ��                >      
 �           �   ��                �   ��                �   ��                �   ��                   ��                
   ��                   ��                   ��                   ��                   ��                %   ��                ,   ��                3   ��                =   ��                D   ��                >       �           M   ��                U      �          [     �          `    t�  �   {       f    ��  �   �       m    ��  �   �      q   ��                >       �           z   ��                >      0 �           C      8 �           H      @ �           �   ��                �    ��  �   _       >      X �           C      ` �           H      p �           �     P �           �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                    ��                >      x �              ��                   ��                   ��                >      � �              ��                >      � �           "   ��                >      � �           #   ��                >      � �              ��                >      � �              ��                >      � �           )   ��                >      � �           1   ��                >      � �           8   ��                >      � �           >   ��                G   ��                >      � �           C      � �           P   ��                >      � �           C      � �                ��                Y    ` �           o    ��  �   T       w    �4  �         �    в  �   \       �    �m  �   �       �    ��  �   {       �    j�  �   9       �    ��  �   ;       �    �  �   �       �    �  �   �       �    �3  �   �       �    |�  �   7      �
    ҳ  �   �       �     �          �    ��  �   �      �    ��  �   �       �    �  �           5    i  �   �       �    �  �           �    Z�  �   P       �    L�  �   �       �    � �              B�  �   �       �    
�  �   �            �              ^  �   �          %�  �   U       !    �y  �   u       /    ��  �   w       6    ��  �   9       ;    � �          A    d�  �   9       G    ��  �   ^       O    ` �          Y    ��  �   �       
    ��  �   �       _    ��  �   [      e    �E  �   :      q    H  �   �       M	    u�  �   �       �    ��  �   w       �    v  �   �       �    
}  �   �      �    h�  �   L       �    '�  �   v      *    ,�  �   �       �    ��  �   U       �    �  �   \       �    T�  �   Y       �    ��  �   M       �    d�  �   K       �      �          �    � �          �    �v  �   �      �    ��  �   <       �    ��  �   �       �    z�  �   L          ��  �   G      
    ( �              K$  �             �8  �   ]      4    �i  �   �       >    ו  �   K       E     �  �           J    }j  �   �      S    (z  �   �      Z       �           c    �"  �   Z      m    �b  �   �       s    �.  �   A       z      �   �       �    ɀ  �   2      �    /-  �   �       �    ��  �   2      �    0 �          �    ��  �   �       �    *'  �   �       �    ��  �   �       �    E�  �   �       �    ��  �   O       �    l�  �   5      �    /  �   i       �    ��  �   P       �
    3�  �   �       �    �-  �   �       �    %�  �   z       �    �6  �   �      N     @ �           �    T�  �   �           ��  �   Y       
    X  �   9           �I  �   �      "     �  �   �      �
    +�  �   9       '    8 �          -     �  �          B	    � �           6    � �          <       �           C    @ �          L     @ �           R    
�  �   �       Y    V3  �   9       c    ~0  �   g       q	    ��  �   D       �    �  �   '       q    �  �   >       w    i�  �   T       ~    �  �   V       �    ��  �   �       �    �/  �   U       �    �g  �         �    Z�  �   n       �    
�  �   }       �    \g  �   �       �    j�  �   �       �    1�  �   9       �    � �          �    o�  �   S       �    'l  �   j      �    	f  �   k       �    ;  �         C	    � �               ��  �   W           Q  �   H          ��  �   �           Ǵ  �   �       &    tf  �   �       2    G  �          =    �_  �          H    ��  �   X       R    n,  �   �       Y    �H  �   �       j    ��  �   ]       p    � �          w    �>  �   D      �    � �          �    �1  �   �      �    ��  �   �       �    ��  �   �       �     �  �           �    �  �   9       �    ��  �   ;       �    �  �   b       �    H �          �    <"  �   �       �    ��  �   K       �    ��  �   *       �    ��  �   K       �    4�  �   �       �	    +�  �   /       �    (  �   r       �     �  �           �    P �          �    S�  �   �       �    ��  �   a       �    \  �         �	    "�  �   S       	    �u  �   +           �*  �   �      	    &  �   �       	    �  �   l       f    �(  �         (	     �  �   �       H	    ��  �   9       /	    jy  �   I       5	    WS  �   e      A	    � �           G	    �  �   9       L	    `�  �   K       �    	�  �         R	    Mn  �         a	    ;�  �   Z       h	    @�  �   6      p	    u�  �   9       u	    ��  �   �       z	    7�  �   2       
    ��  �   �       �	    X �          �	    �M  �   i      �	    ��  �   �       �	    i%  �   �       �	    �X  �   '      �	    J�  �   �       �     �  �           �	    ` �          �	    �  �   S       �	    �&  �   p       �	       �   @      �	    N   �           �	    �c  �   C      �	    ��  �   :       �	    �  �   u      �	    ��  �   �       �	    �  �   ]       �	    h �          M     @ �           
    ��  �   \      
    ��  �   L       
    ��  �   Y       �
       �           
    �`  �   �       '
    ��  �   7       ,
    p �          3
    �W  �   a       =
    ��  �   U       j    �t  �         B
    VX  �   �       �	    (p  �   �      K
    0  �   i       U
    Z�  �   ;       \
    I�  �   3      c
    `   �   �      h
    lo  �   �       y
    v�  �   L       �
       �           �
    ��  �   U       �
    �u  �   9       �
    �0  �   �       �
    
�  �   '       �
       �           �
    x4  �   ^       �	    ��  �   �       �
    ��  �   4       �
    ��  �   a       �
    �  �   �       �
    <�  �   9       �
    �  �   +      �
    ��  �   =       �
    ��  �   �      �
    ��  �   r       �
    k/  �   U       �
    #�  �   L       �
    �a  �   O       lib/setup.asm HEADER_MAGIC HEADER_FLAGS header crt0.c test.c .LC0 .LC1 .LC2 file.c cfs.c alloc_spin_lock pipe.c path.c gui.c font8x16.c window.c bmp.c font.c border.c memcmp.c memcpy.c memset.c strcasecmp.c strcat.c strchr.c strcmp.c strcpy.c strcspn.c string.c strlen.c strncasecmp.c strncmp.c strncpy.c strpbrk.c strrchr.c strsep.c strspn.c strtok.c last.1481 strstr.c strdup.c memmove.c strcoll.c strerror.c ctype.c tolower.c toupper.c stdio.c fopen.c fclose.c fflush.c fputc.c fgetc.c fgets.c fputs.c fread.c fwrite.c remove.c rewind.c fseek.c feof.c ftell.c vfprintf.c vf vsprintf.c vsnprintf.c sn_buf putchar.c sscanf.c perror.c vfscanf.c character _buf.1638 fvalue _buf.1650 ungetc.c getchar.c freopen.c tmpnam.c _tmpnam rename.c itoa.c i2hex.c malloc.c calloc.c free.c realloc.c lldiv.c strtol.c atoi.c atol.c strtoul.c exit.c getenv.c qsort.c qscmp qses qsexc qstexc qs1 system.c strtod.c ftoa.c _precision .LC3 atof.c strtof.c strtold.c abs.c ltoa.c utoa.c srand.c errno.c gmtime.c localtime.c strftime.c clock.c math.c pow.c sqrt.c atan.c acos.c asin.c floor.c ceil.c exp.c locale.c signal.c setjmp.c _GLOBAL_OFFSET_TABLE_ longjmp read_directory_blk drawstring strcpy log sqrt setjmp put clean_blk_enter strtok_r stdout vsprintf ungetc pwd_ptr argv strerror utoa_r __m_i memmove __tm __realloc_r atol __window_puts getenv ceil errno floor strtold _infinity qsort fgets file_update file_read_block memcpy __window_clear BitMAP2 perror ltoa_r tolower system feof malloc remove fs_directory __window_putchar ldexp vsnprintf strtoul itoa __pipe__ stdgetc_r update_directory_entry _drawline fflush argc drawrect BitMAP eh_frame stdputc_r upath tell_r strncasecmp border write_r strtol user rename flush_r strrchr utoa calloc strtod rewind_r atof seek_r strcat read_directory_entry debug_o fseek __free_block_r open_dir ftoa stdin font8x16 __m_c _start obj_list __end strstr write_blk get_file_name atan2 signal strcoll strncmp write_sector draw_char_transparent pow strncpy put_pixel strcasecmp log10 _BLK_ realloc drawchar path_count open_file_r strtok remove_blk memcmp sscanf getfilename file_close pipe_write sigaction read_r file_write_block fread _ctype open_file addr search_blk_null strdup fopen sysgettmpnam localtime memset pwd main ftell srand fclose getchar close_r __data ptr_mouse2 __free_r update_window getkeyw _vsputs_r strcmp color remove_file __bss atan fgetc drawchar_trans strtof strcspn asin ltoa setlocale stderr create_file strsep getkey __malloc_r mouse fputc open_r A__ call_function getpathname strftime i2hex lldiv fwrite __window vfscanf rewind freopen pipe_read exit pipe_r __block_r atoi __heap_r assert_fn gmtime strspn ctr0 drawstring_trans strlen __code toupper wcl filename_cmp clock read_super_block abs strchr fputs acos strchrnul frexp vfprintf strpbrk read_sector free setpath  .symtab .strtab .shstrtab .text .data .got .got.plt .bss .eh_frame .comment                                                                                     �           �                             !              �  �    �                                      '               �         `                              ,             ` �   `                                  5             � �   x     �                             :                �                                         D      0                @     *                                                   0@     �(      	   �                 	                      �h                                                        �s     M                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ELF          >       �   @       `t         @ 8  @  
                 �      �    �       �                    �       �  �    �  �   x        0                            �      �                          Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��  ���_ cole _          �      �            @ �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           I��H�p �   L�H�P �   H�H� �  �   L�H��  �   L�#H��  �   L�+�   �����H��H��H��H��L�������UH��AWSH��@��H�����I���      L�H�}�H�u�H�U�H�M�L�E�L�M�H���������H�H�U�H�H�     H�E�H�H�E�H��     H�H��     H�H� H��H�      H�H��     H�H��H��     H�H��     H�H�@H��H��     H�H�E�H��     H�H�E�H��     H�H�E�H��     H�H�     H�H��H��     H�I�߸    H�yI������H���H��     H�    H���������H�H� H��H��     H�H���������H�H� H��H���������H�H� H�։�I��H��������H��ЉE�E��I��H���������H��АH��@[A_]���UH��AWSH��   ��H�����I��      L�H������Hǅ����    Hǅ����    H�������    �>   H���H�H������H��������H�4H��I��H��������H���H�E�H�}� u�    �}H�U�H������H�Ѻ�  �   H��I��H�͊������H��ЉE�E�H�Ƅ���� H������H��H�
�������H�<I�߸    H���������H��ҁ}��  ~뉐�   H��   [A_]���UH��AWSH�� ��H�����I���      Lۉ}�H�uЃ}�9H�E�H� H��H��������H�<I�߸    H���������H��Ҹ   �   �E�   �   �E�H�H��    H�E�H�H� H��H��������H��Ѓ���tM�E�H�H��    H�E�H�H�H�E�H� H��H� �������H�<I�߸    H���������H��Ѹ   ��E��E�;E��r����    H�� [A_]���UH��AWSH����H�����I���      Lۉ}�H�u�H�E�� ��H�E��@9�sH�E��P#H�E��@9�r"H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@��u)H���������H�H��E�H�։�H�������H���H�E�H�PH�E��@#��H�H�E�H�PH�E�H�@�U�H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  H�E��@��u0H���������H�H� H��t�E�����I��H��g������H��ЋE�H��[A_]���UH��H����H�����I���      L�H�}��E�    H�E�@��u]H�E�@'�PH�E�P'��H�E�P#H�E�@'9�r�H�E�H�PH�E�@'��H��H�H�E�H�PH�E�H�@� ���E��   H�E�@��tH�E�@��uiH�E�@#��u������ZH�E�P'H�E�@#9�r������AH�E�H�PH�E�@'��H�H�E�H�PH�E�H�@� ���E�H�E�@'�PH�E�P'�E�����UH��H����H�����I�h�      L�H���������H�H� H�E��E�    H�E��@��uWH�E��P#H�E��@'9�w�    �AH�E�H�PH�E��@'��H�H�E�H�PH�E�H�@� ���E�H�E��@'�PH�E��P'�E�����UH��H����H�����I���      L�H���������H�H� H�E��E�    H�E��@��uXH�E��@'�PH�E��P'��H�E��P#H�E��@'9�r�H�E�H�PH�E��@'��H��H�H�E�H�PH�E�H�@� ���E��E�����UH��AWH��(��H�����I��      L�H�}�H�u�H�U����u�    �(H�M�H�U�H��H��I��H��/������H���H�E�H�E�H��(A_]���UH��AWSH�� ��H�����I���      L�H�}�H�}� u
������   H�}� tH�E؋@����tH�E��@"<t������zH�E؋@%�   ��u�    �cH�E؋@#H�U؋J�    ��E�H�E؋@��@��u�U�H�E؉�H��I��H�:������H���H�E�H��I��H��6������H��ЉE�E�H�� [A_]���UH��AWSH����H�����I���      L�H�}�H�}� u������0H�E�H��H�M������H���H�E�H��I��H�28������H���H��[A_]���UH��AWSH�� ��H�����I�K�      Lۉ}�H�u�H�}� u
�������  H�EЋ@��u
�    �  H�EЋ@��tH�EЋ@��tH�EЋ@��u!H�UЋE�H�։�H�������H����y  H�EЋ@����unH�EЋP#H�EЋ�+  9�wYH�EЋ�+  ��tKH�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��E�U�H�EЉ�H��I��H�29������H����H�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U܈H�E�� ��H�EЋ@��9�r3H�EЋ@����H�EЉPH�E�f�   H�E�H��H�M������H���H�EЋ@#�PH�EЉP#H�EЋP#H�EЋ�+  9�vH�EЋ�+  �PH�EЉ�+  H�EЋ@���H�EЉP�    H�� [A_]���UH��AWH��(��H�����I�0�      L�H�}�H�}� u
������  H�E؋@��u
�    �v  H�E؋@��tH�E؋@��tH�E؋@��u"H�E�H��H�n������H��ЉE�E��0  H�E؋P#H�E؋�+  9�r
������  H�E؋@����ulH�E؋P#H�E؋�+  9�wWH�E؋�+  ��tIH�E؋@����H�E؉PH�E؋@#H�U؋r�    ���E�U�H�E؉�H��I��H�29������H���H�E؋@#H�U؋J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@� ���E�H�E�� ��H�E؋@��9�rH�E؋@����H�E؉PH�E�f�   H�E؋@#�PH�E؉P#�E�H��(A_]���UH��SH��H��H�����I�b�      L�H�}ȉuĉU�H�M�H�}� u�    �y�E�    H�E�H�E��E�    �FH�E�H��H��������H��ЉE؃}��u�E�    �u��4H�E�H�PH�U��U؈�E��E��E��E��E�9�w��E�    �u�H��H[]���UH��SH��H��H�����I���      L�H�}ȉuĉU�H�M�H�}� u�    �l�E�    H�E�H�E��E�    �9H�E�H�PH�U�� ���E�H�U��E�H�։�H��������H��ЃE��E��E��E��E�9�w��E�    �u�H��H[]���UH��H����H�����I���      L�H�}�H�u��U�}�tZ�}�|�}� t�}�t�nH�E���H�E��P#H�E���H�E��P'�RH�E��@#H�U��H�E��P#H�E��@'H�U��H�E��P'�(H�E���+  H�U�)Љ�H�E��P#H�E��P#H�E��P'�H�E��@#H�U��J�    ��Љ�H�E�f��    ����UH��H����H�����I��      L�H�}�H�}� u�    �	H�E��@#������UH��H����H�����I���      L�H�}�H�}� t7H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@����H�E��P������UH��H��(��H�����I�f�      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H��(��H�����I��      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H����H�����I���      L�H�}��E�_   �(�E�Hc�H�E�H�� < u�E�Hc�H�E�H��  �m��}� y����    ����UH��H����H�����I�S�      L�H�}�H�E�H�E�H�E�H�E��H�E�� </uH�E�H��H�E�H�E�H�E�� ��u�H�E�����UH��H��0  ��H�����I���      L�H������H������H������H�E�H������H�E�H������H�E��E�    �?H�E�� ��u�E�Hc�H�E�H��  �H�E�H�PH�U��U�Hc�H�U�H�� ��E��}�_~��E�    �-H�E�H�PH�U��H�E�H�PH�U�� 8�t�   ��E��}�_~͸    ����UH��SH�� ��H�����I��      L�H�}�H�u�H�E؋PH�E؋@ЉE�E�H�U����H�@     H�H�¾   H�� ������H��ЉE�}� t
�������   �E�    ��   �E�%�  ��H�@     ��H؋���uf�E�%�  ��H�@     ��H��������E�H�U����H�@     H�H�¾   H�� ������H��ЉE�}� t������r�E��m�E�%�  =�  uE�E��E�H�U����H�@     H�H�¾   H�� ������H��ЉE�}� t�������E�H�E؋@$9E����������H�� []���UH��H����H�����I�{�      L؉}��u�H�U�H�M�    ����UH��AWSH��0��H�����I�?�      Lۉ}�H�u�H�U�H�EȋPH�Eȋ@ЉE�H�Eȋ@ �E܉E�ЉE�   �    H�@     H�<I��H�+v������H����E�    �B�U�E�Љ�H�EЋ ��H�@     H��   H�� ������H��ЉE��}� u�E�H�EȋP �E�9�w���H��0[A_]���UH��H����H�����I�Y�      L�H�}�H�u�H�U��R��H�U����H�U�H��H��   I�� ������J� ������UH��AWSH��`��H�����I���      L�H�}�H�u�H�U�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�E�H�E�H�E�H��I��H�,W������H��ЉE�H�E��@,�E��9  H�E�H�E��H�E�� </uH�E��  H�E��H�E�H�E�� ��u׋U�H�E��@ H�M��	��H�M���H�� ������H��ЉE؃}� t#H�E�H��I��H�F�������H��и    ��   �E�    �f�E���Hc�H�E�H�H�E�H�E��@a��t5H�E��@b����@��t#H�E�H�U�H��H��H�"������H��ЉE���E������}� t�E��}�?~����}� u+�}�?%H�EЋ@k�E�H�E��@ �E؉E�ЉE�m��	�E�    �
�}� �����H�E�H��I��H�F�������H��ЋE�H��`[A_]���UH��AWSH��P��H�����I���      L�H�}�H�u�H�U��M�L�E�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�Eغ    �    H��I��H�+v������H��ЋU�H�E��@ H�M��	��H�M؉�H�� ������H��ЉE�}� t#H�E�H��I��H�F�������H��и������   �E�    �T�E���Hc�H�E�H�H�E�H�E��@a��t#H�E�H�U�H��H��H�"������H��ЉE���E������}� t�E��}�?~����}� u:�}�?4�E���Hc�H�E�H�H�EȺ�   H��H��I��H��u������H�����E�����H�E�H��I��H�F�������H��ЋE�H��P[A_]���UH��AWSH��P��H�����I��      L�H�}�H�u�H�U�H�E���C  ��u
������	  H�E���C  ��@v/H�@�������H�<I�߸    H���������H��Ҹ������  H�E��PH�E��@ЉE�H�E���?  H�E��@ �ЋE�ЉE�    I��H���������H���H�E�H�Eغ    �    H��I��H�+v������H��ЋU�H�E��@ H�M��	��H�M؉�H�� ������H��ЉEԃ}� t!H�E�H��I��H�F�������H��ЋE��  H�E���C  ��H��H��H�E�H�H�E�H�EȺ`   �    H��I��H�+v������H���H�E�H��+H��H��!������H���H��H�E�H��H��I��H��x������H����E�    �"H�UȋE�H����uH�UȋE�H�� �E��}�_~�H�E��@` H�E���+  H�EȉPo�U�H�E��@ H�M��	��H�M؉�H�� ������H��ЉE�H�E�H��I��H�F�������H��ЋE�H��P[A_]���UH��AWSH��`��H�����I���      L�H�}�H�u�H�U��S  I��H���������H���H�E�H�EкS  �    H��I��H�+v������H���H�E��PH�E��@ ��H�EЉP�    I��H���������H���H�U�H�BH�E��PoH�EЉ�+  H�E��PH�EЉ�/  H�E��P H�EЉ�3  H�E��H�EЉ�G  �    I��H���������H���H�U�H��K  H�E�H��K  �    �    H��I��H�+v������H���H�E��@k�E�    I��H���������H���H�E��E������E�    �E�    ��  �   I��H���������H���H�U�H��K  �M�Hc�H��H�H�H�E�H��K  �U�Hc�H��H�H� H�E�H�E��   �    H��I��H�+v������H����E�    �<  H�E��@ �E��H�E��@�H�E��P�E�H�H�4�    H�E�H�ʉH�EЋ�;  �PH�EЉ�;  �E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E�;E�ts�E�H�U����H�U�H��H�¾   H�� ������H��ЉE��}� t:H�E�H��I��H�F�������H���H�E�H��H�28������H��и    �   �E��E�H�E��@�����E�    ��U�E�H��    H�E�HЋ �E�}��u	�E�������E��}��  ������}��t�E��}��  � �����H�E�H��I��H�F�������H���H�E�H��`[A_]���UH��AWSH��p  ��H�����I�:�      L�H������H�������   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H������H�E�H��H��I��H��T������H���H�U�H�E�H��H��I��H��W������H��п�   I��H���������H���H�      H�H�      H���   �    H��I��H�+v������H��п   I��H���������H���H�E�H�EȺ   �    H��I��H�+v������H���H�E�H�E�H�E��   �    H��I��H�+v������H����E�    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ ���    Hǅ���    Hǅ���    Hǅ���    Hǅ ���    Hǅ(���    Hǅ0���    Hǅ8���    Hǅ@���    HǅH���    HǅP���    HǅX���    Hǅ`���    Hǅh���    Hǅp���    Hǅx���    H�E�    H�E�    H������H������H��H��I��H��x������H���������<wt������<au�E�   H�E��@   H�E��     H�U�H�E�H��H��H��%������H��ЉE�}� t_H�      H�H��I��H�F�������H���H�E�H��I��H�F�������H���H�E�H��I��H�F�������H��и    �  H�E�H�U�H�M�H�E�H��H��H��%������H��ЉE��}� u_H�      H�H��I��H�F�������H���H�E�H��I��H�F�������H���H�E�H��I��H�F�������H��и    �  H�EȋU��P,H�      H�H�M�H�U�H�u�I�ȹ    H��H�(������H��ЉE�}����   �}� tqH�      H�H������H�U�H�u�A�    H��H��>������H���H�      H�H������H�U�H�u�I�ȹ    H��H�(������H��ЉE�}� ��   H�      H�H��I��H�F�������H���H�E�H��I��H�F�������H���H�E�H��I��H�F�������H��и    ��  �}� t_H�E�H��I��H�F�������H���H�      H�H��I��H�F�������H���H�E�H��I��H�F�������H��и    �r  H�      H�H�U�H�M�H��H��H�5,������H���H�E�H�}� ��   H�      H�H��H�E�H��+�`   H��H��I��H��u������H���H�E�H��+H��H�8!������H���������<wt������<+t������<au
H�E��@"�H�E��@"H�E��@   H�EȋP,H�E���?  H�      H��PsH�E���C  ������<auH�      H��PoH�E��P#H�E�H��I��H�F�������H���H�      H�H��I��H�F�������H���H�E�H��I��H�F�������H���H�E�H��p  [A_]���UH��AWSH��@��H�����I���      L�H�}��   I��H���������H���H�E�H�E�   �    H��I��H�+v������H���H�E�H�E�H�E�   �    H��I��H�+v������H���H�E��@   H�E��     H�U�H�E�H��H��H��%������H��ЉE܃}� t H�E�H��I��H�F�������H��и�����AH�U�H�M�H�E�H��H��H��)������H��ЉE�H�E�H��I��H�F�������H��ЋE�H��@[A_]���UH��AWSH�� ��H�����I���      L�H�}�H�E�H�@H��I��H�F�������H����E�    �TH�E�H��K  �U�Hc�H��H�H� H��t?H�E�H��K  �U�Hc�H��H�H� H��I��H�F�������H��ЃE��}��  ~���H�E�H��K  H��I��H�F�������H���H�E�H��I��H�F�������H���H�E�    �    H�� [A_]���UH��H�� ��L�����I���      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H�� ������I� ������UH��H�� ��L�����I���      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H�� ������I� ������UH��AWSH��   ��H�����I��      L�H��x���H��p�����l����   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H��x���H�E�H��H��I��H��T������H���H�U�H�E�H��H��I��H��W������H��п   I��H���������H���H�E�H�EȺ   �    H��I��H�+v������H���H�E�H�E�H�E��   �    H��I��H�+v������H���H�E��@   H�E��     H�U�H�E�H��H��H��%������H��ЉE��}� t_H�      H�H��I��H�F�������H���H�E�H��I��H�F�������H���H�E�H��I��H�F�������H��и�����-  H�E�H�U�H�M�H�E�H��H��H��%������H��ЉE��}� u_H�      H�H��I��H�F�������H���H�E�H��I��H�F�������H���H�E�H��I��H�F�������H��и�����  H�EȋU��P,H�EȋPH�Eȋ@ЉE�H�EȋP,H�Eȋ@ �ЋE�ЉE��    I��H���������H���H�E�H�E��    �    H��I��H�+v������H��ЋU�H�Eȋ@ H�M��	��H�M���H�� ������H��ЉE��E�    �E�    �   �E���Hc�H�E�H�H�E��E�;�l���}~H�E��@a��ta�E���Hc�H��p���H�H�E���   H��H��I��H��u������H��ЋE���Hc�H��p���H�H��H�8!������H��ЃE����E��}�?�e�����H�E�H��I��H�F�������H���H�E�H��I��H�F�������H���H�E�H��I��H�F�������H��ЋE�H�Đ   [A_]���UH��AWSH��`��H�����I�(�      L�H�}�H�u�H�U�H�M�D�E�H�E�H�E�H�Eغ�   �    H��I��H�+v������H���H�E�H��H��!������H���H��H�E�H��H��I��H��x������H����E�    �"H�U؋E�H����uH�U؋E�H�� �E��}�_~�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉEп    I��H���������H���H�E�H�EȺ    �    H��I��H�+v������H��ЋU�H�E��@ H�M��	��H�Mȉ�H�� ������H��ЉEă}� t!H�E�H��I��H�F�������H��ЋE���  �E�    �$�E���Hc�H�E�H�H�E�H�E��@a��t�E��}�?~���H�E��@a���G  �}�?�=  �U�H�E؉PsH�E��@a��E���H�E؈PbH�U�H�E�H��H��H��"������H���H�U؉BkH�E؋@k���uOH�E�H��H�\�������H�<I�߸    H���������H���H�E�H��I��H�F�������H��и   ��   �E���@��t$H�E؋@kH�U�H�M�H�Ή�H��$������H���H�M�H�E຀   H��H��I��H��u������H��ЋU�H�E��@ H�M��	��H�Mȉ�H�� ������H��ЉEĐH�E�H��I��H�F�������H��и    �JH�E�H��I��H�F�������H���H�E�H��H���������H�<I�߸    H���������H��Ҹ����H��`[A_]���UH��AWSH��P��H�����I���      Lۉ}�H�u�H�U��    I��H���������H���H�E��E�    �E��E��E������E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E��E܋E�;E���   �}� tV�E�H�U����H�U�H��H�¾   H�� ������H��ЉẼ}� t#H�E�H��I��H�F�������H��и�����?  �E�H�U����H�U�H��H�¾   H�� ������H��ЉẼ}� t#H�E�H��I��H�F�������H��и������   �E��E�E��E��E�   H�E��@�����E�    ��U�E�EȋE�H��    H�E�HЋ �E�E�H��    H�E�H��     �}��uL�E�H�U����H�U�H��H�¾   H�� ������H��ЉE̐H�E�H��I��H�F�������H��ЋE��6�E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��Y���H��P[A_]���UH��AWSH��   ��H�����I�t�      L�H��h����   I��H���������H���H�E�H�E�H�E�H�E�H   H�E�H��h���H�E�H��H��I��H��T������H���H�U�H�E�H��H��I��H��W������H��п   I��H���������H���H�E�H�E��   �    H��I��H�+v������H���H��p���H�E�H�E��   �    H��I��H�+v������H���H�E��@   H�E��     H�U�H�E�H��H��H��%������H��ЉE�}� t<H�E�H��I��H�F�������H���H�E�H��I��H�F�������H��и    ��  H�E�H�U�H�M�H�E�H��H��H��%������H��ЉE��}� u<H�E�H��I��H�F�������H���H�E�H��I��H�F�������H��и�����d  H�E��U��P,H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE��    I��H���������H���H�E�H�E��    �    H��I��H�+v������H��ЋU�H�E��@ H�M��	��H�M���H�� ������H��ЉE�}� tSH�E�H��I��H�F�������H���H�E�H��I��H�F�������H���H�E�H��I��H�F�������H��ЋE��l  �E�    �   �E������E���Hc�H�E�H�H�E�H�E��@a��t!H�E�H�U�H��H��H�"������H��ЉE�}� u9H�E��@a �U�H�E��@ H�M��	��H�M���H�� ������H��ЉE�}� ��E��}�?�k����}� tPH�E�H��I��H�F�������H���H�E�H��I��H�F�������H���H�E�H��I��H�F�������H��ЋE��uH�E��@kH�U�H�M�H�Ή�H�2B������H��ЉE�H�E�H��I��H�F�������H���H�E�H��I��H�F�������H���H�E�H��I��H�F�������H��ЋE�H�Đ   [A_]���UH��H����H�5����I��      Lމ}�E�E��}� u�E��   �E����rH�P     H�H�P     H�����UH��H����H�����I���      L�H�}��   H�E�H���r�����UH��AWH����H�����I�y�      L�H�@     H�H�U�H�H     H�    H�        �    H�M�   �    H��I��H�+v������H��ѐH��A_]���UH��AWSH��P��H�����I��      Lۉ}��u��}� u
�    ��  H�H     H�H=�   v%H���������H�<I�߸    H���������H��ҐH�        ���u�H�        ��PH�        ��E����E�E�%�  ��t�E��E�    �E�    �E�    �}� t�E��   �E�   �K  �}��  �=  H�@     H�H�E�H�E�    �E�    �  H�E؋@����   H�E؋@9E���   H�E�H�H�E؋@��H�H�E�H�E؋@+E���H�E؉PH�E؋P�E��H�E؉PH�E�H�E�H�@     H�H�E��E�    �mH�E؋@��tH�E��E��WH�E�H�E�H�E�H�E�H�E�H�@H�PH�E�H�PH�E��@   H�E�H�U�H�H�E��U��PH�E�H�U�H�P�E���!�}��   ~��H�E��E��}��   ������E�   ���}� ��   H�@     H�H�E��E�    �~H�E؋@��tH�E��E��hH�E�H�E��E��H��H������H���H�E�H�E�H�U�H��E��E���H�E��PH�E��U��P�E���+E���H�E��PH�E�H�@   ��}��   �u���H�        �    H�H     H�H�PH�H     H�H�E�H��P[A_]���UH��SH��(��H�����I�̲      L�H�}�H�}� ��  �H�        ���u�H�        ��PH�        �H�E�H�E�H�@     H�H�E��E�    �M  H�E�H� H9E�tH�E��E��2  H�E�H�E�H�H     H�H�P�H�H     H�H�E؋@��uH�E�H��H�@I������H����   H�E؋@��uH�E�H�@H�E�H�E�H�@H�P�H�E�H�PH�E�H�@H��tH�E؋@����   H�E�H�@H��uRH�E�H� H��H�@I������H���H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    ��}��   �������H�        �    ��H��([]���UH��AWH��H��L�����I�ʰ      M�H�}��u�H�E�    �E�    H�}� u�E��   ��H� J������I� ���8  �H�        A� ��u�H�        A� �PH�        A� H�@     I� H�E�H�E�H�E��E�    �   H�E�H� H9E�t
H�E��   H�E�H�E��E�   H�E��P�E��=   v@H�H     I� �U�H�E�H��H��������I�< M�Ǹ    I���������M�A����H�E�H� H�E�H�E��P�E��H�E��P�E��}��   �X���H�        A�     �}� u�E��   ��H� J������I� ���H�E�H��HA_]���UH��H�� ��H�����I�*�      L�H�}�H�u��E�    H�E�H�E��   H�E�� ��H�E��@9�sH�E��P#H�E��@9�rH�E��@#    H�E�f�   H�E�H�PH�E��@#��H�H�E�H�PH�E�H�PH�U�H�U�H�R� �H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  �E��}��E����E�����UH��H�� ��H�����I�*�      L�H�}�H�u��E�    H�E�H�E�H�E��@'�PH�E��P'H�E��P'H�E��@9�rH�E��@'   �H�E��P#H�E��@'9�r�H�E��@'�P�H�E��P'�JH�E�H�PH�E��@'��H�H�E�H�PH�E�H�PH�E�H�HH�M���H�E��@'�PH�E��P'�E��}�~��E�����UH��AWSH��0��H�����I�C�      L�H�}�H���������H�H� H�E�H�E�H�E�H�E�H��I��H��{������H��ЉE�H�E�H��I��H��{������H��ЉE؋U܋E��=   ~
������   H�E�� </uH�E��E�H�HE�H�m�H�E�� </tH�E�H�E�H�PH�U�� /�H�E�H�U�H�E�H��H��I��H��x������H���H�E�H��I��H��{������H��Љ�HE�H�m�H�E�� </u	H�E��  �H�E�H�E��  �    H��0[A_]���UH��AWSH����H�����I���      L�H���������H�H� H��I��H��{������H��Ѓ�w
�    �   H���������H�H� H�E�H�E�H��I��H��{������H��Љ�HE��H�E�H�P�H�U��  H�E�� </u�H���������H�H� H��I��H��{������H��Ѓ�vH�E��  �    H��[A_]���UH��AWSH��0��H�����I��      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
�    ��  H�E�H��I��H��{������H��ЉE�E�H�H�P�H�E�H�� </u�E�H�H�P�H�E�H��  �}� 
�    �  �}���   H�E�H��� <:u%H�U�H�E�H��H��I��H��x������H����K  H�<�������H�<I��H� �������H���H��H�E�H��H��I��H��x������H���H�E�H��I��H��{������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H��x������H����   H�<�������H�<I��H� �������H���H��H�E�H��H��I��H��x������H���H�E�H��I��H��{������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H��x������H���H�E�H��0[A_]���UH��H����H�����I�Ȩ      L�H�}�H�E�H�E�H�}� u�    �+�E�    �H�E�� </u�E�H�E�H�E�� ��u�E�����UH��AWSH��0��H�����I�Z�      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
������   H�E�H��I��H��{������H��ЉE�E�H�HE�H�m��H�E�� </tH�m�H�E�� ��t�E�P��U�����H�E�H�U�H�E�H��H��I��H��x������H���H�E��  �    H��0[A_]���UH��H��0��H�����I�u�      L�H�}�H�u��U܉M�L�E�H���������H�H� H�E��E�H9E�}?H�E��@��H9E�}0H�E�H�E��E�H�E�H��H�E�H�H��    H�E�HE؉������UH��SH��@��H�����I�ަ      Lۉ}ԉuЉỦM�L�E�L�M�f�E�  H�E�H�@H�E�H�E��@�E�}�u�E�    �E�    �   f�E� H�E��@�EȉE��H�H� H�E�H�� f�E�H�E�� ���E��J�E�f#E�f��t5�UЋE��Hc��UԋE��H�H�}��M�U�I��H��H�X������H���f�e�m��}� y��E�H�E��@9E��b�����H��@[]���UH��AWSH��0��H�����I�ǥ      Lۉ}܉u؉UԉM�D�E�L�M��E�    �X�E�    �CH�E�L��   �M�H�E��P�u؋E��Hc��}܋E��H�H��I��H�X������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I��      Lۉ}܉u؉UԉM�D�E�L�M��E�    �p�E�    �[H�E�H��   �E��E�i��E��A��H�E��P�M؋E��Hc��M܋E��H�I��D��H��I��H�X������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I�Q�      Lۉ}܉u؉UԉM�D�E�L�M��}� �[  �}� �Q  �E�    �>H�E�L��   �M�H�E��P�E�Hc��}܋E��H�H��I��H�X������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E����Hc��}܋E��H�H��I��H�X������H��ЃE��E�;E�|��E�    �AH�E�H��   �M�H�E��P�u؋E��Hc��E�H�I��H��I��H�X������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E��Hc��}܋E����H�H��I��H�X������H��ЃE��E�;E�|���H��0[A_]���UH��AWSH��@��H�����I���      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}��  �E�    ��   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��   �E�f#E�f��tDH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�X������H����BH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�X������H���f�e�m��}� �[����E�H�E��@9E��	�����H��@[A_]���UH��SH��8��H�����I�?�      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H�J]������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I���      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}���   �E�    �   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��W�E�f#E�f��tBH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�X������H���f�e�m��}� y��E�H�E��@9E��T�����H��@[A_]���UH��SH��8��H�����I�d�      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H�p_������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I���      L�H�}ȉuĉU��M�D�E�D�M�H���������H�H� H�E�H�E�H   � �? �    H��I��H�+v������H����E�    �U�H�E��P4�UH�E��P8�UH�E��P<H�E��@H   H�E��@L   H�E��P<H�E��PP�UH�E��PTH���������H�H��H�E�H�PXH�E��@D    H�E��PDH�E��P@�U�H�E��P�U�H�E��P�U�H�E��P �U�H�E��P�U H�E��P`�} u�E�   H�E��@�P�H�E��P(H�E��P�E�)ЍP�H�E��P$H�E��@0   �E����H�E��P,H�E��@��H�E��@��H�E�I���Ѻ    �    I��H��q������H���H�E��@4��H�E��@����H�E�I��A�ȹ   �   �   H�*Z������H��Ѓ}� u:H�E��@����H�E�I��A���� �   �   �   H�*Z������H����8H�E��@����H�E�I��A���� �   �   �   H�*Z������H��Ѓ}� t}H�E��@����H�U��E�I��A���� ����   �   H�*Z������H���H�E��@4��H�E��@���ƋE��H�U�I��A�ȹ   ��ƿ   H�*Z������H���H�E��@8A��H�E��@$��H�E��@(��H�E��@,��H�E��@0��H�E�I��H�*Z������H���H�E�H��I��H��{������H������E�H�E�H�pHH�E��@��E܉������)Љ�H�E�H���u�I��A���� ������   ��H��H��`������H���H��H�E��@����H�E�I��A�    �   �   �   H��[������H���H�E�H�PHH�E��@��H���u�I��A���� ������   �ƿX   H�p_������H���H��H�E�H�PHH�E��@��(H���u�I��A���� ������   �ƿ-   H�p_������H���H��H�E�H�e�[A_]���UH��AWSH��0��H�����I�"�      L�H�}�H�u�H�E��P0H�E��@Ѓ�P�E�H�E��P,H�E��@Ѓ��E��E�P   �E�   �E�    �E���� H�E�H��I��H��{������H��ЉE�H�E�L�@H�M؋U܋E���������p��E�<�E��������ƋE���)ƋE��H�E�H���u�M��A�ȉщ�H��H��^������H���H���H�e�[A_]���UH��H����H�����I��      L�H�}��   H�E�H���r�����UH��H����H�����I��      L�H�}������UH��H����H�����I���      L�H�}�H�U��BD    H�U��JDH�U��J@H�U��R8A��H�U��R$��H�U��R(A��H�U��R,��H�U��R0��H�U�I��D��I�*Z������J��А����UH��SH��(��L�����I�,�      Mډ�f�E�H���������I�H� H�E�H���������I�H��H�E�H�PXH�E�@(�P�H�E�@H���к    ��E�H�E�@$�P�H�E�@L���к    ��E�H�E�P<H�E�PPH�E�PD�E�9�rH�E��@D    H�E�@@�PH�E�P@H�E�P@�E�9�r9H�E��@D    H�E�PDH�E�P@H�E�H��H�:g������I����E��  f�}���   H�E�@D����   H�E�@D�P�H�E�PDH�E�H�xHH�E�pTH�E�@PH�U�J,H�U�RLA��H�U�R@A��ʃ���H�U�J0H�U�RHA��H�U�RDA��ʃ�A��H���u�I��A������D�޿    H�J]������I���H����   f�}�	uH�E�@D�PH�E�PD��   f�}�
u!H�E��@D    H�E�@@�PH�E�P@�   f�}���   H�E�H�xHH�E�pTH�E�PPH�E�H,H�E�@LA��H�E�@@A��ȃ���H�E�H0H�E�@HA��H�E�@DA��ȃ�A���E�H���u�I��A���щ�D�މ�H�J]������I���H��H�E�@D�PH�E�PD�E�H�]�����UH��H����H�����I�g�      L؉}�H���������H�H� H�E��U�H�E��P<�����UH��SH��(��H�����I��      L�H�}�H�}� t=H�E�H�E��&H�E�H�PH�U�� f�����H��g������H���H�E�� ��u���H��([]���UH��AWSH��P��H�����I���      L�H�}��u��U��M�L�E�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H�@�������H�<I�߸    H���������H��Ҹ�����6  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H�N�������H�<I�߸    H���������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�f�������H�<I�߸    H���������H��Ҹ   ��   �E�    �   �E�    �   �}� tNH�E�H��   H�E��P�M��E���E��Hc��M��E���E��H��M�I��H��I��H�X������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�X������H��ЃE��}� �U����E��}� �;����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��P��H�����I�đ      L�H�}��u��U��M�D�E�L�M�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H�@�������H�<I�߸    H���������H��Ҹ�����3  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H�N�������H�<I�߸    H���������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�f�������H�<I�߸    H���������H��Ҹ   ��   �E�    �   �E�    �   �}� tKH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�X������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�X������H��ЃE��}� �X����E��}� �>����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��0��H�����I��      Lۉ}܉u؉U�H�M��E�    �   �E�    �t�U�������E��H���������H�Hڋ��E�}� tBH�E�H��   H�EȋP�MԋE��Hc��M؋E��H��M�I��H��I��H�X������H��ЃE��}�~��E��}��o�����H��0[A_]���UH��AWSH��@��H�����I��      Lۉ}̉uȉUĉM�L�E��E���� �E�``` �E���� �EĉE��ẺE܋E��E؋EȉEԋE؍P��E��xH�M��E�I��A�    �   ��I��H��[������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H��[������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H��[������H��ЋEԍP��E܍pH�M��E�I��A�    �Ѻ   ��I��H��[������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H��[������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H��[������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H��[������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H��[������H��ЋEԍP��E܍p�M��E�ȃ�H�M�I��A�    �Ѻ   ��I��H��[������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H��[������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H��[������H��ЋE؍P��M܋E�ȍp��E���H�M�I��A�    �   ��I��H��[������H��АH��@[A_]���UH��H��8��H�����I�֊      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �CH�E�H�PH�U�� ���E�H�E�H�PH�U�� ���E�E�+E�E�}� u�}� t
�m��}� u��E�����UH��H��8��H�����I�@�      L�H�}�H�uЉŰẺE�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M����E��P��U���u�H�E�����UH��H�� ��H�����I�ɉ      L�H�}���U��E�E��E�H�E�H�E��H�E�H�PH�U��U��m��}� u�H�E�����UH��AWSH��0��H�����I�d�      L�H�}�H�u�H�E�H�E�H�E�H�E��E�    H�E�H�PH�U�� ����I��H�̈́������H��ЉE�H�E�H�PH�U�� ����I��H�̈́������H��ЉEԋE�+EԉE܃}� u�}� t뗋E�H��0[A_]���UH��AWSH����H�����I���      L�H�}�H�u�H�E�H��I��H��{������H��Љ�H�E�H�H�E�H��H��I��H��x������H���H�E�H��[A_]���UH��H�� ��H�����I�2�      L�H�}�u�H�E�H�E��H�E�� ��9E�uH�E��H�E�H�E�� ��u۸    ����UH��H�� ��H�����I�ч      L�H�}�H�u�H�E�H�E�H�E�H�E��3H�E��H�E�� 8�u!H�E�� ��H�E�� ��Ѕ�u�    �'H�E�H�PH�U��H�E�H�PH�U�� 8�t����������UH��H��0��H�����I�7�      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E��  H�E�����UH��AWH��(��H�����I���      L�H�}؉uԋU��҉Uԃ}� uOH�U�H��I��H��{������H��҉�H�E�H���   H�E�� ��tH�E�� ��9E�u	H�E��   H�E�H�E؃�H��űE�i��E�H�E�H�E��H�E�H�E� ������H�E� ��!�%������u%H�E� 3E䍐����H�E� 3E���!�%������t�H�E�H�E��H�E�H�E�� ��tH�E�� ��9E�u�H�E�H��(A_]���UH��H��@��H�����I���      L�H�}�H�u�H�U�H�U�H�U������   H�U�H�������   H�E�    H�E�    H�E�    H�E�    �H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�t�H�E�H+E��'H�U����H�Uȉ�H��H�8y������H���H+E�����UH��H����H�����I�[�      L�H�}�H�E�H�E��H�E�H�E�� ��u�H�E�H+E�����UH��AWSH��@��H�����I��      L�H�}�H�u��U�H�E�H�E�H�E�H�E��E�    �kH�E�H�PH�U�� ����I��H�̈́������H��ЉE�H�E�H�PH�U�� ����I��H�̈́������H��ЉEԋE�+EԉE܃}� u�}� t
�m��}� u��E�H��@[A_]���UH��H��(��H�����I�G�      L�H�}�H�u��U�H�E�H�E�H�E�H�E��}� u)������2H�E�H�PH�U��H�E�H�PH�U�� 8�u�m��}� u����E�����UH��H��8��H�����I�ǂ      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �!H�U�H�BH�E�H�E�H�HH�M����E��E�9E�w�H�E��  �E�����UH��AWH����H�����I�H�      L�H�}�H�u�H�M�H�U�H��H��I��H�cz������H��҉�HE�H�E�� ��tH�E���    H��A_]���UH��AWH��(��H�����I�ց      L�H�}؉u�H�U�H��I��H��{������H��҉E��U�H�E�H�H�E��E�    �H�E�� ��9E�uH�E��H�m��E��E�9E�wڸ    H��(A_]���UH��H��0��H�����I�E�      L�H�}�H�u�H�E�H� H�E�H�}� u�    �vH�E�H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u,�}� u
H�E�    �H�E�H���  H�E�H�U�H�H�E���}� u������UH��H��@��H�����I���      L�H�}�H�u�H�E�H�E�H�E�    H�E�    H�E�    H�E�    H�E�� ��u
�    ��   H�E�H��� ��u+�H�E�H�E��H�E�� 8�t�H�E�H+E��   H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�u�H�E�H+E�����UH��H��8��H�����I�U      L�H�}�H�u�H�U�H�}� uH�E�H� H�E�H�}� u
�    ��   �H�E�H�PH�U�� ���E�H�E�H�E��
�E�;E�u��H�E�H�PH�U�� ���E��}� uۃ}� uH�E�H�     �    �   H�E�H��H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u4�}� u
H�E�    �H�E�H��H�E�H�E��  H�E�H�U�H�H�E���}� u������UH��H����H�����I�~      L�H�}�H�u�H�u�H�M�H�(       H�H��H���������H�������UH��AWSH�� ��H�����I��}      L�H�}�H�u�H�E�H��I��H��{������H��ЉE��2�U�H�M�H�E�H��H��I��H�u������H��Ѕ�uH�E��H�E�H�E�� ��uø    H�� [A_]���UH��AWSH�� ��H�����I�,}      L�H�}�H�E�H��I��H��{������H��Ѓ��E�E��I��H���������H���H�E�H�}� u�    �$�U�H�M�H�E�H��H��I��H��u������H��АH�� [A_]���UH��H��8��H�����I��|      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��U�H�E�H�H�E�H�E�H;E�v[H�E�H;E�sQH�E�H�E��E�HE��H�m�H�m�H�E��H�E��H�E�H;E�u��'H�U�H�BH�E�H�E�H�HH�M���H�E�H;E�u�H�E�����UH��AWH����H�����I��{      L�H�}�H�u�H�M�H�U�H��H��I��H�#x������H���H��A_]���UH��AWH����H�����I�u{      Lډ}�H���������H�<I�׸    H���������H�������UH��H����H�����I�'{      L؉}��U���H���������H�Hc��������t�E� �E�����UH��H����H�����I��z      L؉}��U���H���������H�Hc��������t�m� �E�����UH��AWSH��0��H�����I�zz      L�H�}ȉuĉU��M��U�H�E�H��H���������H�<I�߸    I���������I�A��H�E�H��I��H�}�������H���H�E�H�E� �E�H�E� 9E�u��H��0[A_]���UH��AWSH�� ��H�����I��y      L�H�}�H�u�H�E�� ��u�    �LH�E�� <wuH�E�H��I��H���������H���H�U�H�E�H��H��I��H��������H���H�E�H�E�H�� [A_]���UH��AWH����H�����I�Cy      L�H�}�H�U�H��I��H�4������H���H��A_]���UH��AWH����H�����I��x      L�H�}�H�U�H��I��H�M������H���H��A_]���UH��AWH����H�����I��x      L؉}�H�u�H�M��U�H�Ή�I��H��������H���H��A_]���UH��AWSH�� ��H�����I�Yx      L�H�}�H�}� u������VH�E�H��I��H��������H��ЉE�H�E؋@��u+H���������H�H��E�H�։�I��H��������H��ЋE�H�� [A_]���UH��AWH����H�����I��w      L؉}�H�u�H�M��U�H�Ή�I��H�E�������H���H��A_]���UH��AWH����H�����I�ow      L�H�}�H�U�H��I��H���������H���H��A_]���UH��AWSH��@��H�����I�#w      L�H�}ȉu�H�U�H�}� u	H�E��  H�E�H�E�H�E�H�E��E�    H�E�H��I��H��������H��ЉEԃ}����   H�E��@��u7�}�u�}� ~+H���������H�H��E�H�։�I��H��������H��Ѓ}�
tk�E�;E�}E�}�u�}� ~H�E�H;E�vH�m��m��:�}��^���H�E�H�PH�U�UԈ�E��D����}�u�}� ~�m���E��)�������}�~	H�E��  ��Eԉ�H�E�H�E�H��@[A_]���UH��AWSH�� ��H�����I��u      L�H�}�H�u�H�}� u�    �^�E�    �2�E�Hc�H�E�H�� ��H�U�H�։�I��H�E�������H��ЃE�H�E�H��I��H��{������H��ЋU�9�w��E�H�� [A_]���UH��AWH��(��H�����I�%u      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I��������I�A��H��(A_]���UH��AWH��(��H�����I��t      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I�R������I�A��H��(A_]���UH��AWH����H�����I�kt      L�H�}�H�U�H��I��H�zD������H���H��A_]���UH��AWH����H�����I� t      L�H�}�H�U�H��I��H�% ������H��ҐH��A_]���UH��AWH��(��H�����I��s      L�H�}�H�u��U܋U�H�u�H�M�H��I��H�������H���H��(A_]���UH��H����H�����I�}s      L�H�}�H�}� u������!H�E��P#H�E���+  9�r�������    ����UH��AWH����H�����I�"s      L�H�}�H�U�H��I��H��������H���H��A_]���UH��AWSH��`  ��H�����I��r      L�H������H������H�������E�    �E�    �  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H���������H���	E�}���  �E�H��    H��f  H�H��f  H�>��H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E��E�H������H�։�I��H�0�������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�}� t(H������H�E�H��H��I��H�)�������H����O  H������H��H���������H�<I��H�)�������H����   H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E�H�������E�H�։�I��H��������H���H������H������H��H��I��H�)�������H����w  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������
   H��H��I��H�h�������H���H������H������H��H��I��H�)�������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������   H��H��I��H�5�������H���H������H������H��H��I��H�)�������H����  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�EȾ   H��fHn�I��H�#�������H���H������H������H��H��I��H�)�������H����]  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eк
   H��H��I��H���������H���H������H������H��H��I��H�)�������H����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ
   H��H��I��H�h�������H���H������H������H��H��I��H�)�������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ   H��H��I��H�h�������H���H������H������H��H��I��H�)�������H����G  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�E�   H��fHn�I��H�#�������H���H������H������H��H��I��H�)�������H����   H������H�ƿ%   I��H�0�������H��ЋE�Hc�H������H�� ��H������H�։�I��H�0�������H����4�E�Hc�H������H�� ��H������H�։�I��H�0�������H��ЃE��E�Hc�H������H�� ��������    H��`  [A_]���UH��H����H�����I�Hj      L؉��E��E�    �E��S��%wa��H��    H��_  H�H�|_  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��i      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H��������L��Љ�<�����<���H���   A_]���UH��H�� ��H�����I��h      L�H�}�H�u�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E�����UH��AWSH��  ��H�����I�Ah      L�H������H������H��x����E�    H������H�E�f�E�  �E� �E�    �/  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H���������H���	E܃}���  �E�H��    H�^  H�H�^  H�>��H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E��E�H�U�H�E�H��H��H�A�������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H�}� t'H�U�H�E�H��H��H�A�������H���H�E��e  H�E�H���������H�4H��H�A�������H���H�E��7  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E�H�������E�H�։�I��H��������H���H������H�E�H��H��H�A�������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������
   H��H��I��H�h�������H���H������H�E�H��H��H�A�������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������   H��H��I��H�5�������H���H������H�E�H��H��H�A�������H���H�E��3  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�E��   H��fHn�I��H�#�������H���H������H�E�H��H��H�A�������H���H�E��x  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�E��
   H��H��I��H���������H���H������H�E�H��H��H�A�������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ
   H��H��I��H�h�������H���H������H�E�H��H��H�A�������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ   H��H��I��H�h�������H���H������H�E�H��H��H�A�������H���H�E��e  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�Eо   H��fHn�I��H�#�������H���H������H�E�H��H��H�A�������H���H�E��   H�E�H���������H�4H��H�A�������H���H�E�fǅ����  �E�Hc�H������H�� ������H������H�E�H��H��H�A�������H���H�E��8�E�Hc�H������H�� �E�H�U�H�E�H��H��H�A�������H���H�E��E��E�Hc�H������H�� �������H�E��  H�U�H������H)�H��H�Ā  [A_]���UH��H����H�����I�r_      L؉��E��E�    �E��S��%wa��H��    H��V  H�H��V  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��^      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H���������L��Љ�<�����<���Hc�H�����H��  ��<���H���   A_]���UH��AWH���   ��L�����I��]      M�H����������H�����H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H����������H�����H��M��H��������L��Љ�<�����<���H���   A_]���UH��AWSH��0��H�����I��\      L�H�}؉u�H�U�H�M��}�   v
�    �   H�U�H�E�H��H�@       H�<I��H���������H��ЉE�}���  ~�   �I�E�E�}� ~:�U�H�E�H�@       H�4H��I��H��u������H��ЋE�Hc�H�E�H��  �E�H��0[A_]���UH��AWH����H�����I��[      L؉}�H���������H�H�
�U�H�Ή�I��H�E�������H���H��A_]���UH��AWSH�� ��H�����I��[      L�H�}�H�}� tj�E�    �?H���������H�H��E�Hc�H�E�H�� ��H�։�I��H�E�������H��ЃE�H�E�H��I��H��{������H��ЋU�9�w���H�� [A_]���UH��AWH���   ��L�����I��Z      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H��������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I�Z      M�H��8���H��0���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�H���������I�<M�׸    H���������L�������UH��AWH����H�����I�gY      L�H�}�H�U�H��I��H�O�������H��ҐH��A_]���UH��AWH��(��H�����I�Y      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H�Έ������H��Ѹ    H��(A_]���UH��AWH��(��H�����I��X      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H�Έ������H����H�E�H�E�� < tH�E�H   H9E�sH�E�� <
u�H�E��  H�E�H;E�����H��(A_]���UH��AWSH��0��H�����I�X      L�H�}�H�uЉỦM�H�@      H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H�Έ������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H�@      H�H�E�H�@      �0H�@      �D �}�u-�U�H�E�    H��I��H���������H���H�U�H��   �}�u+�U�H�E�    H��I��H���������H��Љ�H�EЉ�[�}�u,�U�H�E�    H��I��H���������H��Љ�H�E�f��)�U�H�E�    H��I��H���������H��Љ�H�EЈ�    H��0[A_]���UH��AWSH��0��H�����I�oV      L�H�}�H�uЉỦM�H�@     H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H�Έ������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H�@     H�H�E�H�@     �0H�@     �D �}�u'H�E�H��I��H��������H����Z�H�E�� �+�}�u%H�E�H��I��H��������H���fH~�H�U�H��    H��0[A_]���UH��SH��8��H�����I�4U      L�H�}�H�u�H�U��E�    �E�    ��  �E�    �E�Hc�H�E�H�� ������%��  �E��E�Hc�H�E�H�� ������lu�E��E�   �E�Hc�H�E�H�� ����H��������H���	E�}��o  �E�H��    H�1M  H�H�&M  H�>��H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H�צ������H�����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H�<�������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�ާ������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�ާ������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H����?  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�ާ������H�����   H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�ާ������H����jH�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H���������H������E��E�Hc�H�E�H�� ��������E�H��8[]���UH��H����H�����I��P      L؉��E��E�    �E��S��%wa��H��    H� J  H�H�J  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I�*P      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I�?O      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��H����H�����I�ON      L؉}�H�u�H�}� u������w�}��u������jH�E��@#��tH�E��@#�P�H�E��P#H�E��@#H�U��J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U���E�����UH��AWSH����H�����I��M      L�H���������H�H� H��I��H��������H��ЉE�}��t+H���������H�H��E�H�։�I��H��������H��ЋE�H��[A_]���UH��AWH��(��H�����I�M      L�H�}�H�u�H�U�H���������H�<I�ϸ    H���������H�������UH��H����H�����I��L      L�H�}��	   H�E�H���r�����UH��SH����H�����I�}L      L�H�}�H�}� u.H�@     H�<H�=�������H���H�@     H��H�E�H��H�=�������H���H�E�H��[]���UH��AWSH��0��H�����I��K      L�H�}�H�u�H�E�H���������H�4H��I��H��������H���H�E�H�}� u
������   �E�    H�E�H��I��H��{������H��ЉE܃}�`~	�E�   �$H�E�H�P+H�E�H��H��I��H��x������H���H�E��@���H�E��PH�E�H��I��H���������H��ЋE�H��0[A_]���UH��H��0��H�����I�K      L؉}�H�u�H�E�H�E��E܉E��E�    �}� y,H�E�H�PH�U�� -�}�   �u�E�����E���E��؉E�H�E�H�E�M�Hc�Hi�gfffH�� ��������)�����)��ʉЍH0H�E�H�PH�U�ʈ�E�Hc�Hi�gfffH�� ����)ЉE�}� u��}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWSH��@��H�����I��I      L�H�}�H�u��U�H�}� u#H�E�H�E�H�E�H�PH�U�� 0H�E��  �  H�E�H�E؋E�Hc�H�E�H�H�E��3H�E؃��E�H�m��}�	~�7   ��0   �U��H�m���H�E�H�E�H;E�wËE�Hc�H�E�H��  H�E�H�E��E�    �8H�E�� <0uH�E��"H�U�H�E�H��H��I��H��x������H�����E��E�;E�|�H�E�H�E�H�E�H��I��H��{������H��Љ�H�E؋E�H�U�)Љ�H�M�H�E�HȾ    H��I��H�+v������H���H��@[A_]���UH��AWH����H�����I�HH      L؉}�U�    ��I��H� J������H���H��A_]���UH��AWH����H�����I��G      L؉}�u�U��U��I��H���������H���H��A_]���UH��AWH����H�����I��G      L�H�}�H�U�H��I��H�'M������H��ҐH��A_]���UH��AWH����H�����I�`G      L�H�}�u�M�H�U��H��I��H�(O������H���H��A_]���UH��H����H�����I�G      L؉}�u�E��}�E��E��}�ЉE��}� x�E���y�E����E��E�+E�E��!�}� y�E���~�E����E��U��E�ЉE�H�E�����UH��H�� ��H�����I��F      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H�� ��H�����I��E      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H��H��H�����I�3E      L�H�}�H�u��U�H�E�H�E�H�E�H�PH�U�� ���E�E���H���������H�H������ ��uǃ}�-u�E�   H�E�H�PH�U�� ���E��"�E�    �}�+uH�E�H�PH�U�� ���E�}� t�}�u9�}�0u3H�E�� <xtH�E�� <XuH�E�H��� ���E�H�E��E�   �}� u�}�0u�   ��
   �E��}� t	H��   ������H�E�E�Hc�H�E�H�H��H�ЉE؋E�Hc�H�E�H�H��H�E�}� t�}� ~�E�)E�H�E��]�H�E�    �E�    �E���H���������H�H��������t�m�0�[�E���H���������H�H���������5  �E���H���������H�H��������t�7   ��W   )E�E�;E���   �}� ��   �}� tgH�E�H;E�|H�E�H;E�u0�E�;E�~(�E�����H�E�   �H���������H�� �����   �E�   �E�H�H�U�H��H�E��E�H�H)E��eH�E�H;E�H�E�H;E�u-�E�;E�~%�E�����H�E����H���������H�� �����$�E�   �E�H�H�U�H��H�E��E�H�HE���H�E�H�PH�U�� ���E��y������H�}� t�}� t
H�E�H���H�E�H�U�H�H�E�����UH��AWH����H�����I��A      L�H�}�H�M�
   �    H��I��H���������H���H��A_]���UH��AWH����H�����I��A      L�H�}�H�M�
   �    H��I��H���������H���H��A_]���UH��AWAVAUATSH����H�����I�NA      L�H�}�H�uȉU�L�eп    L��L�`� �؉���H���������H�H������ ��uЃ�-u�   L��L�`� �����+uL��L�`� �؃}� t�}�u-��0u(A�$<xt	A�$<XuI�D$� ��I���E�   �}� u��0u�   ��
   �EċE�Hc������    H��I�ǋE�Hc������    H��H�Љ�A�    A�    ����H���������H�H��������t��0�T����H���������H�H��������tz����H���������H�H��������t�7   ��W   )�;]�}GE��x
M9�wM9�u��9�~A������A�   �E�H�L��Hc�I�L��L�`� ���;������E��yA�����H���������H�� "   �	����tI��H�}� tE��tI�D$��H�E�H�U�H�L��H��[A\A]A^A_]���UH��H����H�����I�?      L؉}��   �   ���r����UH��AWSH����H�����I��>      L�H�}�H�E�H���������H�4H��I��H�#x������H��Ѕ�uH���������H�H� ��    H��[A_]���UH��AUATSH�� ��H�����I�X>      L�H�}�H�u�H��     ��E�L�e�H�]�E�,$L��L�`��H��H�XD�(�m��}� uې�H�� [A\A]]���UH��H��8��H�����I��=      L�H�}�H�u�H�U�H��     ��E�H�E�H�E�H�E�H�E�H�E�H�E�H�E�� ���E�H�E�H�PH�U�H�U���H�E�H�PH�U�H�U���H�E�H�PH�U��U���m��}� u�������UH��SH��H��H�����I�3=      L�H�}�H�u�H��     ��E�H�E�H+E��EȋE�9E���  �E�����EȺ    ��E��EȋU�H�E�H�H�E�H�E�H�E�H�E�H�E�E�H�H��H��H�E�H�H�E�H�E�H;E�sjH��     H�H�U�H�E�H��H���щEă}� u/�E�H�H��HE�H�U�H�E�H��H��H���������H�����  �}� y�E�H�HE���  �H�E�H;E���   H��     H�H�U�H�E�H��H���щEă}� u)�E�H�HE�H�U�H�E�H��H��H���������H���뢃}� ��   H�E�H;E�uA�E�H�HE�H�U�H�M�H�E�H��H��H��������H��ЋE�H�HE�H�E�H�E��M���H�U�H�E�H��H��H���������H��ЋE�H�H��HE��E�H�HE���   �E�H�H��HE�����H�E�H;E���   H�E�H+E�H��H�E�H+E�H9�|4�E�Hc�H�E�H�H�E�H��H��H���������H���H�E�H�E������H�U�H�E�H��H��H���������H��ЋE�Hc�H�E�H�H�E������E�H�H��HE�H�U�H�M�H�E�H��H��H��������H��ЋE�H�H��HE�H�E�H�E������H��H[]���UH��H�� ��H�����I�B:      L�H�}��u�U�H�M�H��     H�U�H��U�H��     ��U��U���H�U�H�H�U�H��H��H���������H��А����UH��AWH����H�����I��9      L�H�}�H���������H�<I�׸    H���������H��Ѹ����H��A_]���UH��H��@��H�����I�e9      L�H�}�H�u�H�U�H�U��H�E�H�U����H���������H�Hc���҃� ��u��E�    H�U���҃�+t��-u�E�   H�E�H�����������E��E�    �E�    �E�    �;�M�H�����������Y�H�U���҃�0�*��X��E�H�E��E�H�U����H���������H�Hc���҃���u�H�U����.uuH�E��?�M�H�����������Y�H�U���҃�0�*��X��E�H�E��E��E�H�U����H���������H�Hc���҃���u��U�)U�}� uH���������f���  �}� t�E�H� �������f(fW��E�H�U����etH�U����E��   �E�    H�E�H�U���҃�+t��-u�E�   H�E��E�    �%�M܉����҉�H�U���҃�0ʉU�H�E�H�U����H���������H�Hc���҃���u��}� t�U�)U���U�U�}����|	�}�   ~H� ���������   H�����������E��E�E܃}� yF�]��A�E܃���t&�}� y�E��^E��E���E��YE��E��}��E��Y��E��}� u�H�}� tH�E�H�U�H��E�����UH��H����H�����I�06      L؉}�H�E�   �E�    �H�U�H��H��H�H�H�E��E��E�;E�|�H�E�����UH��AWSH��@��H�����I��5      L��E�H�}��u�H�}� u	H�E��  H�E�H�E�H��������f��f/E�v,H�E�H�PH�U�� -�E�H� �������f(fW��E��E�H�0�������f/s�E��H,�H�E��/�E�H�0���������\��H,�H�E�H�       �H1E�H�E�H�E�H�E�H��x�H*��H��H���H	��H*��X��M��\�f(��EȋE���H���������H���H��x�H*��H��H���H	��H*��X��YE�H�0�������f/s�H,�H�E��*H�0���������\��H,�H�E�H�       �H1E�H�E�H�E�H�M�H�U�H�E�H��������H�43H��I�߸    I�,�������I�A��H�E�H��@[A_]���UH��AWH����H�����I��3      L�H�}�H�U�    H��I��H���������H���H��A_]���UH��AWH����H�����I��3      L�H�}�H�u�H�M�H�U�H��H��I��H���������H����Z�H��A_]���UH��AWH��(��H�����I�:3      L�H�}�H�u�H�M�H�U�H��H��I��H���������H����E��E�H��(A_]���UH��H����H�����I��2      L؉}��E����3E�)�����UH��H��@��H�����I��2      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�    H�}� y>H�E�H�PH�U�� -H�       �H9E�uH��������H�E�H�E��H�E�H��H�E�H�E�H�E�H�M�H�gfffffffH��H��H��H��H��?H)�H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U��ʈH�M�H�gfffffffH��H��H��H��H��?H)�H��H�E�H�}� u�H�}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U߈H�E�H;E�w�H�E�����UH��AWH��8��H�����I�21      L�H�}�H�uЉU�H�U�H�U�H�}� yH�U�H�JH�M��-H�]�H�U�H�U��}�u$H�M�H�u�   H��I��H�5�������H����H�M�H�U�H��H��H�J�������H���H�E�H��8A_]���UH��H��0��H�����I��0      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E�H�M�H���������H��H��H��H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U�ʈH�E�H���������H��H��H��H�E�H�}� u�H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWH��8��H�����I��/      L�H�}�H�uЉU�H�U�H�U�H�U�H�U��}�u$H�u�H�M�   H��I��H�5�������H����H�M�H�U�H��H��H�o�������H���H�E�H��8A_]���UH��H����H�����I��.      L؉}������UH����H�����I��.      Lظ   ]���UH��H����H�����I��.      L�H�}��    ����UH��H����H�����I�w.      L�H�}�H���������H�H� ����UH��H����H�����I�<.      L�H�}�H���������H�H� ����UH��H�� ��H�����I�.      L�H�}��u�H�U�H�M�    ����UH����H�����I��-      Lظ    ]���UH��H����H�����I��-      L��E�H�8�������f������UH��H����H�����I�g-      L��E�H�8�������f������UH��H����H�����I�.-      L��E��}�H�8�������f������UH��H����H�����I��,      L��E�H�}�H�8�������f������UH��H����H�����I��,      L��E��M�H�8�������f������UH��H��(��H�����I�w,      L��E��M��E��U��U��E��E��E������������������������������]��E�����UH��H����H�����I�	,      L��E����E����]��E�����UH��H����H�����I��+      L��E�H�@�������f������UH��H����H�����I��+      L��E�H�H�������f������UH��H����H�����I�\+      L��E�H�P�������f������UH��H����H�����I�#+      L��E�H�X���������E��E�����UH��H����H�����I��*      L��E�H�`�������f������UH��H����H�����I��*      L��E�H�h�������f������UH��H����H�����I�m*      L��E�H�p�������f������UH��H����H�����I�4*      L��E�H�x�������f������UH��AWH����H�����I��)      L��E��E�H���������H�f(�fHn�I��H�}�������H���H��A_]���UH��H����H�����I��)      L؉}�H�u�    ����UH��AWH����H�����I�f)      Lډ}�H�u�H���������H�<I�׸    H���������H�������UH��AWH��(��H�����I�)      Lى}�H�u�H�U�H���������H�<I�ϸ    H���������H�������UH��AWSH�� ��H�����I��(      L�H�}�H���������H�<I�߸    H���������H����E�    �.�E�H�H��    H�E�HЋ ��I��H��������H��ЃE��}�?~̸����H�� [A_]���UH��AWH����H�����I�(      L�H�}�u�H���������H�<I�׸    H���������H�����f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�                                                                          ~ � � � � � � � � ~             ~ � � � � � � � � ~                 l � � � � | 8                   8 | � | 8                   < < � � �   <                < ~ � � ~   <                      < <              � � � � � � � � � � � � � � � �           < f B B f <           � � � � � � � � � � � � � � � �        2 x � � � � x             < f f f f <  ~               ? 3 ? 0 0 0 0 p � �              c  c c c c g � � �               � < � < �             � � � � � � � � � � �               > � >                  < ~    ~ <                f f f f f f f   f f              � � � {                | � ` 8 l � � l 8  � |                       � � � �              < ~    ~ <  ~              < ~                           ~ <                      �                         0 ` � ` 0                         � � � �                       ( l � l (                      8 8 | | � �                   � � | | 8 8                                                 < < <                  f f f $                             l l � l l l � l l           | � � � |   � � |               � �   0 ` � �             8 l l 8 v � � � � v           0 0 0 `                             0 0 0 0 0 0               0         0                   f < � < f                         ~                                    0                     �                                                           0 ` � �             8 l � � � � � � l 8              8 x       ~             | �    0 ` � � �             | �   <    � |               < l � �                 � � � � �    � |             8 ` � � � � � � � |             � �     0 0 0 0             | � � � | � � � � |             | � � � ~     x                                                       0                  0 ` 0                      ~     ~                     ` 0      0 `             | � �                       | � � � � � � � |              8 l � � � � � � �             � f f f | f f f f �             < f � � � � � � f <             � l f f f f f f l �             � f b h x h ` b f �             � f b h x h ` ` ` �             < f � � � � � � f :             � � � � � � � � � �             <         <                   � � � x             � f f l x x l f f �             � ` ` ` ` ` ` b f �             � � � � � � � � � �             � � � � � � � � � �             | � � � � � � � � |             � f f f | ` ` ` ` �             | � � � � � � � � |           � f f f | l f f f �             | � � ` 8   � � |             ~ ~ Z       <             � � � � � � � � � |             � � � � � � � l 8              � � � � � � � � � l             � � l | 8 8 | l � �             f f f f <     <             � � �   0 ` � � �             < 0 0 0 0 0 0 0 0 <               � � � p 8                 <         <          8 l �                                                   �       0                                     x  | � � � v             � ` ` x l f f f f |                   | � � � � � |                < l � � � � v                   | � � � � � |              6 2 0 x 0 0 0 0 x                   v � � � � � |  � x       � ` ` l v f f f f �                 8      <                        f f <       � ` ` f l x x l f �             8         <                   � � � � � � �                   � f f f f f f                   | � � � � � |                   � f f f f f | ` ` �             v � � � � � |                � v f ` ` ` �                   | � ` 8  � |              0 0 � 0 0 0 0 6                    � � � � � � v                   � � � � � l 8                   � � � � � � l                   � l 8 8 8 l �                   � � � � � � ~   �             � �  0 ` � �                 p                                        p         p                       v �                        8 l � � � �                               ��� ��� ~~~                                 uuu ��� ��� ���                                 ��� ��� ��� ��� ;;;                          ��� ��� ~~~ ��� ���                         ��� ��� ���     ��� ���                         ��� ���      ��� ��� ppp                 @@@ ��� ���         III ��� ���                 ��� ��� ��� ��� ��� ��� ��� ���                 ��� ���                 zzz ��� ���         ``` ��� ���                     ��� ���         ��� ��� MMM                     ��� ��� bbb     ��� ���                         ||| ��� ���      ��Cr %s usage: %s FILE...
 %s: failed to open '%s'
        Entrada maior que o limite
 Erro ao criar o arquivo "%s"
       Error ao criar o arquivo "%s", atingio o limite de arquivos na entrada de directorio
   Panic: __malloc, sem espaco na tabela de alocacao
      panic: realoc sem espaco, %lx size = %d %d
 PWD BitMAP error
 Not suport BitMAP 4-bit Not suport BitMAP > 8-bit strerrorr
                      (((((�AAAAAABBBBBB                                �Dubug: %s %x %x
        (null)  1�������[�������ߙ��������������E�������������������������������1�������1�������1�������1�������1�������1�������1�������1�������1�������1�������1�������_��������������Þ������u�������u���������������ɠ������ɠ������ɠ������ɠ��������������ɠ������ɠ������ɠ������ɠ������ɠ������ɠ������ɠ������ɠ������ɠ������ɠ����������������������ɠ����������������������ɠ��������������ɠ������ɠ������ɠ������ɠ������ɠ������ɠ������ɠ������ɠ������ɠ��������������ɠ��������������ɠ������ɠ��������������(null) %        ը���������������������H����������������������L�������L�������ը������ը������ը������ը������ը������ը������ը������ը������ը������ը������ը���������������������i���������������������i�������������������������������������������������������������������������������������������������������������������������������`�������r���������������������������������������r�������������������������������������������������������������������������������i���������������{�������������������������������panic: sscanf()
        ,��������������E����������������������,�����������������������,�������,�������,�������,�������,�������,�������,�������,�������,�������,�������,��������������Z�������,�������õ������õ��������������0�������0�������0�������0��������������0�������0�������0�������0�������0�������0�������0�������0�������0�������0���������������������0�������'��������������0��������������0�������0�������0�������0�������0�������0�������0�������0�������0���������������0��������������0�������0��������������panic: freopen()
 r+ PWD call system funtion error. 
                 $@       �        %lu.%lu                �              �C                                                                        �_�
�@panic: signal()
 panic: sigaction()
 panic: setjmp()  panic: longjmp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �   �  �   �  �   � �    �   � �    �  �   8 �    �  �     �   H �   h �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          zR x�  ,      @ ���   E�CG����B�A�       (   L   ���#   E�CJ���B�A�   (   x   ���   E�CG���B�A�   (   �   ���Z   E�CG��G�B�A�      �   ���   E�C�   �   ����    E�C��      ����    E�C��     0  	��p    E�CF�`�A�$   T  U���    E�CG����B�A�$   |  ��r    E�CG��_�B�A�(   �  ^��   E�CG��	�B�A�   $   �  N
���   E�CF���A�       �  ����    E�CE���A�      ����    E�CE���A�   @  "���    E�C��    `  ���A    E�Cx�      �  ��i    E�C`�        �  F��U    E�CL�    �  {��U    E�CL�    �  ���i    E�C`�      ���g    E�C^�    $  @���    E�C�� $   D  ���   E�CE�{�A�      l  i��9    E�Cp�  $   �  ����    E�CG����B�A�   �  C��^    E�CU� (   �  ���   E�CG���B�A�   (      j���   E�CG����B�A�   (   ,  ��]   E�CG��J�B�A�   (   X  9��   E�CG��l�B�A�   (   �  ���D   E�CJ��.�B�A�   (   �  �"��:   E�CG��'�B�A�   $   �  �#��    E�CG����B�A�     �$���    E�C��    $  >%���    E�C�� (   D  �%���   E�CJ����B�A�   (   p  �)��i   E�CG��V�B�A�   (   �  �,��H   E�CG��5�B�A�   (   �  /��e   E�CJ��O�B�A�      �  G3��a    E�CX�      �3��9    E�Cp�      4  �3���    E�CF�w�A�(   X  4��'   E�CG���B�A�   $   �  �6��   E�CE���A�   $   �  �8���   E�CF���A�      �  R:��    E�C��    �  2;���    E�C�� (     �;��O   E�CG��<�B�A�   $   @  =���    E�CG����B�A�(   h  �=��C   E�CG��0�B�A�      �  �?��k    E�Cb� $   �  ?@���    E�CG����B�A�   �  �@���    E�C�� $   �  uA��   E�CE��A�   $   $  bB���    E�CG����B�A�$   L  �B���    E�CG����B�A�(   t  �C���   E�CG����B�A�   (   �  E��j   E�CG��W�B�A�       �  DF���    E�CE���� (   �  �F��   E�CG���B�A�       	  �G���    E�CE���� (   @	  gH���   E�CG��q�B�A�   $   l	  �L��   E�CG����B�A�   �	  �M��9    E�Cp�     �	  �M��+    E�Cb�     �	  �M���    E�C��     �	  /N���   E�CE����   
  �P��I    E�C@�     8
  �P��u    E�CE�f�A�(   \
  KQ���   E�CG����B�A�   (   �
  T���   E�CG����B�A�   $   �
  �V���    E�CG����B�A�,   �
  lW��2   E�CG���B�A�            nZ���    E�C��    ,  �Z��w    E�Cn�    L  ;[��b    E�CY� $   l  }[���    E�CG����B�A�$   �  \��z    E�CG��g�B�A�   �  b\��a    E�CX�    �  �\���    E�C��    �  ]��{    E�Cr� $     x]��+   E�CF��A�      D  {^��6   E�C-�   d  �_��L    E�CC� $   �  �_���    E�CG����B�A�   �  ]`���    E�Cw�    �  �`��}    E�Ct� $   �  a��r    E�CF�b�A�    $     da���    E�CF���A�       <  �a���    E�C��    \  lb��3   E�C*�   |  c��7   E�C.�   �  �d��W    E�CN� $   �  �d���    E�CG����B�A�$   �  =e���    E�CG����B�A�     �e���    E�C�� $   ,  Wf��V    E�CF�F�A�       T  �f��P    E�CF�       t  �f��U    E�CL�    �  �f��U    E�CL� $   �  g���    E�CG����B�A�$   �  �g���    E�CG����B�A�$     h��K    E�CF�{�A�     $   ,  *h��K    E�CF�{�A�     $   T  Mh��S    E�CF�C�A�    $   |  xh���    E�CG����B�A�$   �  �h��S    E�CF�C�A�    $   �  i��K    E�CF�{�A�     ,   �  6i��[   E�CG��H�B�A�       $   $  aj���    E�CG����B�A�$   L  �j��]    E�CF�M�A�    $   t  k��]    E�CF�M�A�    $   �  Gk��K    E�CF�{�A�     $   �  jk��L    E�CF�|�A�     $   �  �k��Y    E�CF�I�A�         �k��Y    E�CP� $   4  �k��K    E�CF�{�A�     (   \  l���   E�CJ��{�B�A�       �  �t���    E�C��     $   �  u���    E�CI���A�       �  �u��l    E�Cc� (   �  v���   E�CJ����B�A�          �~���    E�C��     $   D  D��   E�CI���A�    $   l  ����    E�CI���A�    $   �  ����    E�CG����B�A�$   �  ����\    E�CF�L�A�    $   �  ǁ���    E�CG����B�A�$     E����    E�CI���A�       4  ����    E�CI�    $   T  ����L    E�CF�|�A�         |  ����e    E�CF�U�A�    �  �����    E�CF���A�(   �  v����   E�CG����B�A�   (   �  ���=   E�CG��*�B�A�   $     ����\   E�CE�M�A�      D  3����    E�C�� $   d  �����    E�CI���A�    $   �  �����    E�CI���A�       �  M����    E�C�� $   �  ߍ���    E�CG��z�B�A�   �  D���Y    E�CF�         }���9    E�Cp�  $   <  �����    E�CE�q�A�    $   d  ����    E�CG����B�A�   �  ����G   E�C>�,   �  ���u   E�CG��b�B�A�       $   �  *���M    E�CF�}�A�     $     O���O    E�CF��A�     $   ,  v���L    E�CF�|�A�     $   T  ����S    E�CF�C�A�       |  Œ���    E�C�    �  -����    E�C��    �  �����    E�C��    �  A���2   E�C)�$   �  S���U    E�CF�E�A�    $   $  ����U    E�CF�E�A�    4   L  ����L   E�CM�����-�B�B�B�B�A�      �  ����7    E�C       $   �  ؙ��w    E�CG��d�B�A�(   �  '���{    E�CI���d�B�B�A�   �  v����    E�C�� $     ����   E�CE���A�       @  Ν���    E�Cx�     $   d  +���\    E�CF�L�A�       �  _���5   E�C,�   �  t���_    E�CV� ,   �  �����   E�CG����B�A�       $   �  n���P    E�CF�@�A�    $   $  ����Z    E�CF�J�A�    $   L  ȣ��^    E�CF�N�A�       t  ����4    E�Ck�     �  ���v   E�Cm�$   �  h����    E�CF���A�       �  ����    E�C�� $   �  Ȧ���    E�CF���A�       $  5���*    E�Ca�     D  ?���'    E�C^�     d  F���/    E�Cf�     �  U���;    E�Cr�     �  p���;    E�Cr�     �  ����:    E�Cq�     �  ����'    E�C^�       ����9    E�Cp�     $  ŧ��9    E�Cp�     D  ާ��<    E�Cs�     d  ����=    E�Ct�     �  ���>    E�Cu�     �  5���n    E�Ce�    �  ����;    E�Cr�     �  ����9    E�Cp�       ����9    E�Cp�     $  Ш��9    E�Cp�     D  ���D    E�C{�     d  ���9    E�Cp�     �  &���9    E�Cp�     �  ?���9    E�Cp�     �  X���9    E�Cp�  $   �  q���a    E�CF�Q�A�         ����2    E�Ci�     ,  ����T    E�CF�   H  ����X    E�CF�$   d  0����    E�CG����B�A�   �  ����T    E�CF�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            GCC: (Ubuntu 9.3.0-17ubuntu1~20.04) 9.3.0                                        �                  �  �                   �                 ` �                 � �                    �                                     ��                     ��_ cole _             ��                )        �           6         �           0    ��                �    ��                7      h �           <      j �           A      m �           F      � �           K    ��                R    ��                7      � �           <      � �           A      � �           �   ��                X     � �          7      8 �           <      p �           h    ��                o    ��                7      � �           v    ��                |    ��                �    ��                �    ��                7      � �           <      � �           A      � �           �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                �    ��                   ��                   ��                   ��                &   ��                0   ��                :   ��                D   ��                M   ��                V   ��                _    � �          i   ��                r   ��                {   ��                �   ��                �   ��                7      � �           �   ��                �   ��                �   ��                �   ��                7        �           �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                    ��                	   ��                   ��                   ��                #   ��                *   ��                2   ��                =    �  �   �       7       �           3   ��                @   ��                =    �  �   �       7       �           <       �           A   ��                L   ��                K   ��                W    � �          ^   ��                �   ��                4   ��                h   ��                7      	 �           q   ��                z   ��                �    7�  �   e       N    ��  �   �       �    >�  �   �      �    � �          �    �  �   =      �    � �          =    {�  �   �       {   ��                |   ��                �   ��                �   ��                �   ��                7       �           �   ��                �    � �   `       �   ��                7      * �           �   ��                �   ��                �   ��                �   ��                   ��                   ��                   ��                   ��                   ��                   ��                #   ��                *   ��                1   ��                ;   ��                B   ��                7      - �           K   ��                S      �          Y     �          ^    ��  �   {       d    r�  �   �       k     �  �   �      o   ��                7      1 �           x   ��                7      P �           <      X �           A      ` �           �   ��                �    $�  �   _       7      x �           <      � �           A      � �           F      p �           �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                7      � �               ��                   ��                   ��                7      � �              ��                7      � �              ��                7      � �              ��                7      � �              ��                7      � �              ��                7      � �           "   ��                7      � �           *   ��                7      � �           1   ��                7      � �           7   ��                @   ��                7      � �           <      � �           I   ��                7       �           <       �                ��                R    ` �           h    3�  �   T       p    Y6  �         �    S�  �   \       �    o  �   �       �    �  �   {       �    ��  �   9       �    K�  �   ;       �    ��  �   �       �    p�  �   �       �    5  �   �       �    ��  �   7      �
    U�  �   �       �     �          �    �  �   �      �    �  �   �       �    �  �           .    �j  �   �       �    �  �           �    ݔ  �   P       �    ��  �   �       �    � �          �    œ  �   �       �    ��  �   �            �          	    �_  �   �          ��  �   U           6{  �   u       (    ��  �   w       /     �  �   9       4    � �          :    ��  �   9       @    �  �   ^       H    ` �          R    �  �   �        
    %�  �   �       X    .�  �   [      ^    XG  �   :      j    �I  �   �       F	    ��  �   �       z    �  �   w       �    <"  �   #      �    �w  �   �       �    �~  �   �      �    �  �   L       �    ��  �   v      #    ��  �   �       �    -�  �   U       �    ��  �   \       �    ל  �   Y       �    
�  �   M       �    �  �   K       �      �          �    � �          �    'x  �   �      �    &�  �   <       �    z�  �   �       �    ��  �   L      �    N�  �   G          ( �              �%  �             8:  �   ]      -    9k  �   �       7    Z�  �   K       >     �  �           C     l  �   �      L    �{  �   �      S       �           \    t$  �   Z      f    ]d  �   �       l    D0  �   A       s    E�  �   �           L�  �   2      �    �.  �   �       �    !�  �   2      �    0 �          �    V�  �   �       �    �(  �   �       �    |�  �   �       �    ��  �   �       �    W�  �   O       �    ��  �   5      �    �0  �   i       �    n�  �   P       �
    ��  �   �       �    f/  �   �       �    ��  �   z       �    n8  �   �      G     @ �           �    ו  �   �       �    ~�  �   Y           �Y  �   9           :K  �   �          ��  �   �      �
    ��  �   9            8 �          &     �  �          ;	    � �           /    � �          5       �           <    @ �          E     @ �           K    ��  �   �       R    �4  �   9       \    2  �   g       j	    1�  �   D       �    ��  �   '       j    ��  �   >       p    ��  �   T       w    ��  �   V           �  �   �       �    C1  �   U       �    ui  �         �    ��  �   n       �    ��  �   }       �    �h  �   �       �    �  �   �       �    ��  �   9       �    � �          �    ��  �   S       �    �m  �   j      �    �g  �   k       �    �<  �         <	    � �           �    6�  �   W           �R  �   H          ~�  �   �           J�  �   �           �g  �   �       +    �H  �          6    *a  �          A    @�  �   X       K    �-  �   �       R    fJ  �   �       c    -�  �   ]       i      �          p    @  �   D      z    � �              O3  �   �      �    %�  �   �       �    y�  �   �       �     �  �           �    ��  �   9       �    �  �   ;       �    ��  �   b       �    H �          �    _#  �         �    0�  �   K       �    ]�  �   *       �    �  �   K       �    ��  �   �       �	    ��  �   /       �    �)  �   r       �     �  �           �    P �          �    ��  �   �       �    Y�  �   a       �    �]  �         �	    ��  �   S       	    ow  �   +           ",  �   �      	    �'  �   �       	    ��  �   l       _    *  �         !	    ��  �   �       A	    u�  �   9       (	    �z  �   I       .	    �T  �   e      :	    � �           @	    ��  �   9       E	    �  �   K       �    ��  �         K	    �o  �         Z	    ��  �   Z       a	    Ê  �   6      i	    ��  �   9       n	     �  �   �       s	    ��  �   2       
    �  �   �       }	    X �          �	    )O  �   i      �	    �  �   �       �	    �&  �   �       �	    `Z  �   '      �	    ��  �   �       �     �  �           �	    ` �          �	    ��  �   S       �	    =(  �   p       �	       �   @      �	    N   �           �	    Ie  �   C      �	    S�  �   :       �	    ��  �   u      �	    w�  �   �       �	    ��  �   ]       �	    h �          F     @ �           �	    �  �   \      
    2�  �   L       
    D�  �   Y       {
       �           
    *b  �   �        
    I�  �   7       %
    p �          ,
    ?Y  �   a       6
    S�  �   U       c    /v  �         ;
    �Y  �   �       �	    �q  �   �      D
    �1  �   i       N
    ��  �   ;       U
    ̏  �   3      \
    `   �   �      a
    �p  �   �       r
    ��  �   L       y
       �           �
    ��  �   U       �
    6w  �   9       �
    h2  �   �       �
    ��  �   '       z
       �           �
    �5  �   ^       �	    E�  �   �       �
    v�  �   4       �
    "�  �   a       �
    ��  �   �       �
    ��  �   9       �
    ��  �   +      �
    b�  �   =       �
    {�  �   �      �
    
�  �   r       �
    �0  �   U       �
    ��  �   L       �
    c  �   O       lib/setup.asm HEADER_MAGIC HEADER_FLAGS header crt0.c .LC0 .LC1 .LC2 .LC3 file.c cfs.c alloc_spin_lock pipe.c path.c gui.c font8x16.c window.c bmp.c font.c border.c memcmp.c memcpy.c memset.c strcasecmp.c strcat.c strchr.c strcmp.c strcpy.c strcspn.c string.c strlen.c strncasecmp.c strncmp.c strncpy.c strpbrk.c strrchr.c strsep.c strspn.c strtok.c last.1481 strstr.c strdup.c memmove.c strcoll.c strerror.c ctype.c tolower.c toupper.c stdio.c fopen.c fclose.c fflush.c fputc.c fgetc.c fgets.c fputs.c fread.c fwrite.c remove.c rewind.c fseek.c feof.c ftell.c vfprintf.c vf vsprintf.c vsnprintf.c sn_buf putchar.c sscanf.c perror.c vfscanf.c character _buf.1638 fvalue _buf.1650 ungetc.c getchar.c freopen.c tmpnam.c _tmpnam rename.c itoa.c i2hex.c malloc.c calloc.c free.c realloc.c lldiv.c strtol.c atoi.c atol.c strtoul.c exit.c getenv.c qsort.c qscmp qses qsexc qstexc qs1 system.c strtod.c ftoa.c _precision atof.c strtof.c strtold.c abs.c ltoa.c utoa.c srand.c errno.c gmtime.c localtime.c strftime.c clock.c math.c pow.c sqrt.c atan.c acos.c asin.c floor.c ceil.c exp.c locale.c signal.c setjmp.c _GLOBAL_OFFSET_TABLE_ longjmp read_directory_blk drawstring strcpy log sqrt setjmp put clean_blk_enter strtok_r stdout vsprintf ungetc pwd_ptr argv strerror utoa_r __m_i memmove __tm __realloc_r atol __window_puts getenv ceil errno floor strtold _infinity qsort fgets file_update file_read_block memcpy __window_clear BitMAP2 perror ltoa_r tolower system feof malloc remove fs_directory __window_putchar ldexp vsnprintf strtoul itoa __pipe__ stdgetc_r update_directory_entry _drawline fflush argc drawrect BitMAP eh_frame stdputc_r upath tell_r strncasecmp border write_r strtol user rename flush_r strrchr utoa calloc strtod rewind_r atof seek_r strcat read_directory_entry debug_o fseek __free_block_r open_dir ftoa stdin font8x16 __m_c _start obj_list __end strstr write_blk get_file_name atan2 signal strcoll strncmp write_sector draw_char_transparent pow strncpy put_pixel strcasecmp log10 _BLK_ realloc drawchar path_count open_file_r strtok remove_blk memcmp sscanf getfilename file_close pipe_write sigaction read_r file_write_block fread _ctype open_file addr search_blk_null strdup fopen sysgettmpnam localtime memset pwd main ftell srand fclose getchar close_r __data ptr_mouse2 __free_r update_window getkeyw _vsputs_r strcmp color remove_file __bss atan fgetc drawchar_trans strtof strcspn asin ltoa setlocale stderr create_file strsep getkey __malloc_r mouse fputc open_r A__ call_function getpathname strftime i2hex lldiv fwrite __window vfscanf rewind freopen pipe_read exit pipe_r __block_r atoi __heap_r assert_fn gmtime strspn ctr0 drawstring_trans strlen __code toupper wcl filename_cmp clock read_super_block abs strchr fputs acos strchrnul frexp vfprintf strpbrk read_sector free setpath  .symtab .strtab .shstrtab .text .data .got .got.plt .bss .eh_frame .comment                                                                                    �           �                             !              �  �    �                                      '               �         `                              ,             ` �   `                                  5             � �   x     �                             :                �                                         D      0                @     *                                                   0@     �(      	   �                 	                      i                                                         t     M                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ELF          >       �   @                  @ 8  @                   �      �    �      �                   �      � �    � �    �       `                   `        �      �    @       @             Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��  ���_ cole _          �      �            ` �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           I��H�P� �   L�H�0� �   H�H� � �   L�H�� �   L�#H�� �   L�+�   �����H��H��H��H��L�������UH��AWSH��@��H�����I�Y�     L�H�}�H�u�H�U�H�M�L�E�L�M�H�P�������H�H�U�H�H���     H�E�H�H�E�H�H�     H�H�H�     H�H� H��H�x�     H�H�h�     H�H��H�8�     H�H�H�     H�H�@H��H�0�     H�H�E�H�P�     H�H�E�H�(�     H�H�E�H�p�     H�H���     H�H��H�@�     H�I�߸    H��������H���H�X�     H�    H�@�������H�H� H��H�`�     H�H�H�������H�H� H��H���������H�H� H�։�I��H�/�������H��ЉE�E��I��H�&�������H��АH��@[A_]���UH��AWH��(��H�����I�~�     L�H�}�H�u�H�UЋ��u&H�E��@�,���H�E؋H�к    ����   H�UЋ��uQH�E�H�@H�E��E�    �,�e�H�E�� ��E�E�H�U؋J�    ��ЉE�H�E�H�E�� ��uɋE��%H���������H�<I��H��!������H��Ҹ����H��(A_]���UH��AWSH��0��H�����I���     L�H�}�H�uЉU�H�E�    H�EЋ ��uqH�E�    H�E�H�@�U�Hc�H��H�H� H�E��?H�E� ��u H�E��@H�E��H.�z	.���   H�E�H�E�H�E�H�@ H�E�H�}� u��   H�EЋ ��u~H�E�    H�E�H�@�U�Hc�H��H�H� H�E��KH�E� ��u,H�E�H�PH�E�H�@H��H��I��H�`E������H��Ѕ�t H�E�H�E�H�E�H�@ H�E�H�}� u�����H�}� u�    �H�E�H��0[A_]���UH��AWSH�� ��H�����I�;�     L�H�}��-H�E�H�@ H�E�H�E�H��I��H���������H���H�E�H�E�H�}� u̐�H�� [A_]���UH��AWSH�� ��H�����I���     Lۉ}ܿ   I��H��������H���H�E�H�}� u'H���������H�<I��H��������H��и    �mH�E�U܉PH�E��  �Eܾ   ��I��H�4�������H���H�U�H�BH�E�H�@H��u'H���������H�<I��H��������H��и    �H�E�H�� [A_]���UH��AWSH�� ��H�����I���     L�H�}��E�    �/H�E�H�@�U�Hc�H��H�H� H��H��������H��ЃE�H�E؋P�E�9�w�H�E�H�@H��I��H���������H���H�E�H��I��H���������H��АH�� [A_]���UH��AWSH�� ��H�����I�5�     L�H�}�H�u�H�U�H�E�H��H��H�t������H��ЉE�}� y
�    ��   �U�H�M�H�E�H��H��H�\������H���H�E�H�}� ��   �(   I��H��������H���H�E�H�}� u'H���������H�<I��H��������H��и    �eH�M�H�E�H�PH� H�H�QH�E��@   H�E�H�@�U�Hc�H��H�H�H�E�H�P H�E�H�@�U�Hc�H��H�H�E�H�H�E�H��H�� [A_]���UH��AWSH�� ��H�����I���     L�H�}�H�E�� �E�    �kH�E�H�@�U�Hc�H��H�H� H�E��BH�E�H��I��H�t������H���H�E�H��H��I��H�t������H���H�E�H�@ H�E�H�}� u��E�H�E؋P�E�9�w���H�� [A_]���UH��AWSH�� ��H�����I�/�     L�H�}؉u�H�E؋P�E�9���   �EԉE��   H�E�H�@�U�Hc�H��H�H� H����   H�E�H�@�U�Hc�H��H�H� �@��t`H�E�H�@�U�Hc�H��H�H� H��I��H��d������H���H�E�H�@�U�Hc�H��H�H� H��H��I��H��d������H����:�E�H�E؋P�E�9��I���I��H�a������H���I��H�a������H���H�� [A_]���UH��AWSH��0��H�����I� �     Lۿ   I��H��\������H���H�Eؿ   I��H��\������H���H�E�H�}� tH�}� u%H���������H�<I��H��������H����u  �   I��H��\������H���H��t%H� �������H�<I��H��������H����4  H�E؋ ��t%H�H�������H�<I��H��������H����  H�E�H�@H�E�H�EЋ ��u!H�EȾ    H��H��������H�����  H�U�H�E�H��H��H�t������H��ЉEă}� ��  H�E�H�@�U�Hc�H��H�H� H�E��N  H�E�H�Mк   H��H��I��H�[B������H��Ѕ��  H�E�H�@ H��u$�EčPH�Eȉ�H��H��������H����"  H�E�H�@ �@��tCH�E�H�@ H��I��H��d������H���H�E�H�@ H��H��I��H��d������H�����   H�E�H�@ H�@ H�E��H�E�H�@ H�E�H�}� tH�E��@��t�H�}� u!�EčPH�Eȉ�H��H��������H����vH�E�H��I��H��d������H���H�E�H��H��I��H��d������H����>H�E�H�@ H�E�H�}� �����H�}� u H���������H�<I��H��������H���H��0[A_]���UH��H����H�����I���     L�H�}�H�PD      H�U�H������UH��AWH����H�����I���     L�H�@D      H�H��I��H��U������H��҉E�}��t�E���    H��A_]���UH��AWH����H�����I�R�     L؉}�H�@D      H��U�H�Ή�I��H��~������H��ҐH��A_]���UH����H�����I���     L�H�HD      H�H�JH�HD      H�H�HD      H�H��� ��]���UH��H����H�����I���     L؉}�H�HD      H�H�J�H�HD      H������UH��AWSH����H�����I�S�     L�H�}�H���     �   H�<������H�<I��H��$������H���H��������H�<I��H�/%������H���H�E�H���������H�4H��I��H�VS������H���H�@D      H�H�@D      H�H��u�   �)H�E�H��I��H�Py������H��Ѕ�t�   ��    H��[A_]���UH��AWS��H�����I�Z�     L�H�@D      H�H��t5H�@D      H�H��I��H��S������H���H�@D      H�    �[A_]���UH��AWSH��P��H�����I���     L�H�}�H���     �   H��������H�<I��H��$������H���H�T������H�<I��H�/%������H���H�HD      H�E�H�H�U�H�E�H���������H�4H��I�߸    H�in������H���H�E�H��I��H�Py������H��Ѕ�t�   ��    H��P[A_]���UH��AWH����H�����I���     L�H�}�H�PD      H�H��tH�PD      H�H�E�H�����>H���������H�H� H�U�H���������H�41H��I�ϸ    I��c������I�A�АH��A_]���UH��H����H�����I�[�     L؉}��u�H�8D      ���~%H���������H�<H��������H��и   �sH�8D      �H�8C      Hc�H�4�M���H�8D      �H�8C      Hc�H��H�H�H�J�U��H�8D      ��JH�8D      ��    ����UH����H�����I���     L�H�8D      ��J�H�8D      ��]���UH��AWAVAUATSH��(  ��H�����I�9�     L�H������H������H������H��H��I��H��E������H���H���     �����  H�8D      ����  H�8D      ���H�8C      H�Hڋ�H���������H�Hc�L�4�H�p�������H�H�H�8D      ���H�8C      H�H��H�H�H��� Hc�H��H�H�H��H�L�(H���     D�$H�������    H��I��H��D������H���M��L��D��H���������H�43H��I�߸    I�in������I�A��H�������    H��I��H��D������H���H�)�������H�4H��I�߸    H�in������H���H�8D      ����E���   H�8C      �E�H�Hڋ�H���������H�Hc�L�,�H�p�������H�H�H�8C      �E�H�H��H�H�H��� Hc�H��H�H�H��H�L� H�������    H��I��H��D������H���L��L��H�@�������H�43H��I�߸    I�in������I�A�Ѓm��}� �2����sI��H�Vz������H���I��H���     D�$H�������    H��I��H��D������H���L��D��H�`�������H�43H��I�߸    I�in������I�A��H������H��H��������H��АH��(  [A\A]A^A_]���UH��H����H�����I��     L�H�}�H��D      H�U�H������UH��H����H�����I���     L�H�}�H��D      H�U�H������UH����H�����I���     L�H�ؾ     H�]���UH��AWSH����H�����I�U�     L��  ����E����#�o  ��H��    H��� H�H��� H�>��I�߸    H�X�������H��҅��g  �    �  H���������H��    �  �f  H���������H��     �  �H  H���������H�� �PH���������H����  �  �  �  �  �  �  �  ��  �  ��  �  ��  �  ��  �  ��  �	  ��  H���������H�� �P�H���������H�f��  �  �
  �  �  �  �  �z  �  �p  �  �f  �  �\  �  �R  �  �H  �  �>  �  �4  �  �*  H�ؾ     H�<I��H��o������H��Љ�H���������H�f��  ��   H�ؾ     H�<I��H�K�������H����Z�H���������H�� �  �   H�ؾ     H�<I��H��m������H��Љ�H���������H�f��  �sH�ؾ     ����`H���     H��U�H���������H�4H��I�߸    H��c������H��Ѹ    H��(������H��҉E�}� �"����    H��[A_]���UH��AWAVAUATSH��8��H�����I�7�     L��E�   H���     ���uH�ؾ     H�H�E��6H���     �    H���     �Hc�H�ؾ     H�H�H�E�H���     L�4H��
      L�,H� �     L�,H�����������
uI��M�e H�ز������H�I9�u7�}� u1I�EH�E�H�}� ��  H�E�H�H�ز������H�H9��q  H��D      H��ЉE�H�E�H�PH�U��U���E�    L�e�L����H�ز������H�9���   �E�H�H� H�E�L�$H��
      H�I9���  A�$H��H��H�H�H��H��H�       H�H�I9��y  A�D$H��H��H�H�H��H��u&H��D      H�H�m�H�E�� �������  A�D$H��H��H�H�H��H��H�       H�L�,L��L�pL�(�D  L����H�ز������H�9���  H�ز������H�L)�H��H�ز������H�H�H�E�L�e��E�H�H�I�H��
      H�I9���   A�$H��H��H�H�H��H��H�       H�H�I9�u}A�D$H��H��H�H�H��H��u&H��D      H�H�m�H�E�� �������u  A�D$H��H��H�H�H��H��H�       H�L�,L��L�pL�(�.  H�8��������E�H�H��H��H� H�E�L�$H��
      H�I9���   A�$H��H��H�H�H��H��H�       H�H�I9�uzA�D$H��H��H�H�H��H��u&H��D      H�H�m�H�E�� �������   A�D$H��H��H�H�H��H��H�       H�L�,L��L�pL�(�HM�mM��tM�e H�ز������H�I9�t�����H��D      H�H�m�H�E�� ��������G������  ��  H�E�H�P�H�U��  I�H����  I�H�@H���     H�H���     H�H���Z  H���     H�� ���B  H���     L�4H���     H�� H�XD      H�H����tw�(I��H��D      H�H�E�H�H�H�M�� ������H���     H�� �؉�I�H�@��H�Ǹ    H�0������H��҃�tH���     H�I9�w�H�E�� ��H���������H���     L�4H�ؾ     H�H�U�H)�H�Ѓ���H���     �H���     �H�ؾ     H�H�� H���     H�H�PH���     H�� �	  H��D      H�H�E�� ������L��L�p�H���     H�H9��%���H�ؾ     ���u&H��
      H��     H�H��    �   H��D      H��Љ�H�ؾ     �H�ؾ     ���H���������H�����������~2H���     H�H���������H�։�I��H��T������H���H�ؾ     H�H�E��Q���H��8[A\A]A^A_]���UH��H����H�����I���     L�H�}��u�H�}� u!�    �)H�E�H�PH�U�� 9E�u�   �H�E�� ��uܸ    ����UH����H�����I���     L�H��D      H���]���UH��AWH����H�����I�[�     L؉}�H���     H��U�H�Ή�I��H��T������H��ҐH��A_]���UH��H����H�����I��     L؉}�H��D      H��E����Ґ����UH��AWATSH��(��H�����I���     L�H�}�H�u�H�E�H��I��H��H������H���A��H�E�H��I��H��H������H���D����   ��I��H�4�������H���H�E�H�}� u'H���������H�<I��H��������H��и    �NH�E�H�PH�U��  H�U�H�E�H��H��I��H��E������H���H��H�E�H��H��I��H��D������H���H��([A\A_]���UH��AWSH�� ��H�����I���     L�H�}�H�E�H��I��H��H������H��Ѓ��   ��I��H�4�������H���H�E�H�}� u'H���������H�<I��H��������H��и    �/H�E�H�PH�U��  H�U�H�E�H��H��I��H��E������H���H�� [A_]���UH��AWSH�� ��H�����I���     L�H�}�H�E؋ ��t'H���������H�<I��H��!������H��и   �rH�E�H�@H�U�H��H��I��H�̓������H����Z�H�E��@H�E�� ��t'H��������H�<I��H��!������H��и   �H�E��    �    H�� [A_]���UH��AWSH�� ��H�����I��     L�H�}�H�E؋ ��u.H��T      H�E�H�PH� H�H�TH��T      H��~H��T      �   H�E؋ ��uTH�E�H�@H�U�H��H��I��H�̓������H����Z�H��T      �DH�E�� ��uH��T      �   H��T      H�H�� [A_]���UH��AWSH����H�����I�$�     L�H�}�H�E� ��t*H�0�������H�<I��H��!������H��и   �  H�E��@�,��*�H�E��H.�zI.�uDH�E��@�,���H�X�������H�4H��T      H�<I�߸    H�in������H����@H�E��@�Z�H�[�������H�4H��T      H�<I�߸   H�in������H���H��T      H�<H�@2������H���H��I��H��w������H���H�U�H�BH�E�H�@H��u�   �H�E��    �    H��[A_]���UH��AWATSH��  ��H�����I���     L�H������H������H�PH������� ����?�c"  ��H��    H�W� H�H�L� H�>��H��
      H�H�PH��
      H��    �h"  H��
      H��    H��
      H�H�PH��
      H�H�����������@�"  H��
      H��    H��
      H�H�PH��
      H�H�����������@��!  H��
      H��    H��
      H�H�PH��
      H�H�����������@�!  H��
      H��    H������H�PH�������H��
      H�H�PH��
      H�3���*��@�'!  H��
      H��    H�������H��
      H�H�PH��
      H�3���*��@H��������   H��
      H��    H��
      H�H�PH��
      H�H��������@H�������   H������� ��������H������H��
      H��    H���������H�H� ������Hc�H��H�H��
      H�H�PH��
      H�3H�H�P�   H��
      H�H��
      H�H�QH��
      H�3H�PH� H�H�Q��  H��
      H�H��
      H�H�QH��
      H�3H�PH�@H�H�Q�  H��
      H�H��
      H�H�QH��
      H�3H�P(H�@ H�H�Q�=  H��
      H�H��
      H�H�QH��
      H�3H�P8H�@0H�H�Q��  H��
      H�H��
      H�H�QH��
      H�3H�PHH�@@H�H�Q�  H��
      H�H��
      H�H�QH��
      H�3H�PXH�@PH�H�Q�w  H��
      H�H��
      H�H�QH��
      H�3H�PhH�@`H�H�Q�5  H��
      H�H��
      H�H�QH��
      H�3H�PxH�@pH�H�Q��  H��
      H�H��
      H�H�QH��
      H�3H���   H���   H�H�Q�  H��
      H�H��
      H�H�QH��
      H�3H���   H���   H�H�Q�c  H��
      H�H������H�PH������� ��H��H�H��
      H�H�AH��
      H�3H�H�RH�H�Q�  H�p�������H�H�H������� ��H��H�H�H��H�H��
      H�H�AH��
      H�3H�BH�RH�H�QH�������  H��
      H�H�P�H��
      H�H��
      H�H��� ��t*H�`�������H�<I��H��!������H��и   �9  H��
      H�H��
      H�H��H�@H��H��I��H��������H���H������H������ u
�   ��  H��
      H�H�H�H������H�PH� H�H�Q�  H��
      H�H�PH��
      H��     �  H��
      H�H��
      H�H�P�H�@�H�H�QH��
      H�H�PH��
      H��6  H��
      H�H�P�H��
      H�H��
      H�H��
      H�H�PH� H�H�Q��  H��
      H�H�P�H��
      H�H��
      H�H��
      H�H�JH�PH� H�H�Q�  H��
      H�H�P�H��
      H�H��
      H�H��
      H�H�J H�PH� H�H�Q�A  H��
      H�H�P�H��
      H�H��
      H�H��
      H�H�J0H�PH� H�H�Q��  H��
      H�H�P�H��
      H�H��
      H�H��
      H�H�J@H�PH� H�H�Q�  H��
      H�H�P�H��
      H�H��
      H�H��
      H�H�JPH�PH� H�H�Q�H  H��
      H�H�P�H��
      H�H��
      H�H��
      H�H�J`H�PH� H�H�Q��  H��
      H�H�P�H��
      H�H��
      H�H��
      H�H�JpH�PH� H�H�Q�  H��
      H�H�P�H��
      H�H��
      H�H��
      H�H���   H�PH� H�H�Q�L  H��
      H�H�P�H��
      H�H��
      H�H��
      H�H���   H�PH� H�H�Q��  H��
      H�H�P�H��
      H�H��
      H�H��
      H�4H������H�HH������� ��H��H�H�H�RH�H�Q�  H��
      H�H�P�H��
      H�H��
      H�H�p�������H�H�0H������� ��H��H�H�H��H�H�H�QH�FH�VH�������  H��
      H�H��0� ��t*H�`�������H�<I��H��!������H��и   ��  H��
      H�H�P�H��
      H�H��0H�@H��H��I��H��������H���H�� ���H�� ��� u
�   �v  H��
      H�H�� ���H�P�H�@�H�H�QH��
      H�H�P�H��
      H��(  H������H�PH������� �������H��
      H������Hc�H��H������H)�H��HЋ ��t*H�`�������H�<I��H��!������H��и   �  H��
      H������Hc�H��H������H)�H��H�H��
      H������Hc�H��H������H)�H��H�H�@H��H��I��H��������H���H�����H����� u
�   �&  H��
      H�H�����H�P�H�@�H�H�QH��
      H�H�P�H��
      H���  H��
      H�H��0� ��t*H���������H�<I��H��������H��и   �  H��
      L�$H��
      H�H�P�H��
      H�H��0H�@H��H��I��H��������H���H��I�D$�I�T$�H�H�QH��
      H�H�P�H��
      H��  H��
      H�H������H�PH������� ��H��H�H�����H��
      H�H9������  �&H��
      H�H�PH��
      H��    H��
      H�H9����w�H��
      H�����H��A  H��
      H�H��� ��u+H��
      H�H��H�����������@�   H��
      H�H��� ��t3H��
      H�H��H��H�
3������H��Ѕ�t
�   ��  H��
      H�H���HH���������f��/�r&H��
      H�H��H�����������@H��
      H�H���@�H,���I��H�"������H���H��
      H�L�b�H��I��H�ix������H���I�D$H��
      H�H��H�@H��u
�   �
  H��
      H�H���    ��  H��
      H�H�� H��(���H��
      H�H��H�� ���H��
      H�H�P�H��
      H�H��(����H�� ���� 9�tH��
      H�H���    ��  H��(���� ����  ��H��    H�� H�H�� H�>��H��
      H�H���    �  H��(����@H�� ����H.�z.�u�   ��   H��
      H�H����[  H��(���H�PH�� ���H�@H9�u�   ��   H��
      H�H����  H��(���H�PH�� ���H�@H9�u�   ��   H��
      H�H�����   H��(���H�PH�� ���H�@H9�u�   ��   H��
      H�H����   H��(���H�PH�� ���H�@H9�u�   ��   H��
      H�H����^H�� ���H�PH��(���H�@H��H��I��H�`E������H��Ѕ�u�   ��   H��
      H�H����
�   �u  H��
      H�H��H�����������@�E  H��
      H�H�� H��8���H��
      H�H��H��0���H��
      H�H�P�H��
      H�H��8���� ��uPH��0���� ��uBH��8����HH��0����@/�v�   ��   H��
      H�H����   H��8���� ��tH��8���H��H��4������H��Ѕ�u,H��0���� ��t(H��0���H��H��4������H��Ѕ�t
�   �8  H��0���H�PH��8���H�@H��H��I��H�`E������H��Ѕ�y�   ��   H��
      H�H���H��
      H�H��H�����������@�  H��
      H�H�� H��H���H��
      H�H��H��@���H��
      H�H�P�H��
      H�H��H���� ��uPH��@���� ��uBH��H����HH��@����@/�r�   ��   H��
      H�H����   H��H���� ��tH��H���H��H��4������H��Ѕ�u,H��@���� ��t(H��@���H��H��4������H��Ѕ�t
�   �  H��@���H�PH��H���H�@H��H��I��H�`E������H��Ѕ��   ��   H��
      H�H���H��
      H�H��H�����������@�'  H��
      H�H�� H��X���H��
      H�H��H��P���H��P���� ��tH��P���H��H�
3������H��Ѕ�u,H��X���� ��t(H��X���H��H�
3������H��Ѕ�t
�   �  H��X����HH��P����@�X�H��X����@H��
      H�H�P�H��
      H��F  H��
      H�H�� H��h���H��
      H�H��H��`���H��`���� ��tH��`���H��H�
3������H��Ѕ�u,H��h���� ��t(H��h���H��H�
3������H��Ѕ�t
�   �
  H��h����@H��`����H�\�H��h����@H��
      H�H�P�H��
      H��e
  H��
      H�H�� H��x���H��
      H�H��H��p���H��p���� ��tH��p���H��H�
3������H��Ѕ�u,H��x���� ��t(H��x���H��H�
3������H��Ѕ�t
�   ��	  H��x����HH��p����@�Y�H��x����@H��
      H�H�P�H��
      H��	  H��
      H�H�� H�E�H��
      H�H��H�E�H�E�� ��tH�E�H��H�
3������H��Ѕ�u&H�E�� ��t%H�E�H��H�
3������H��Ѕ�t
�   �	  H�E��@H�E��H�^�H�E��@H��
      H�H�P�H��
      H��  H��
      H�H�� H�E�H��
      H�H��H�E�H�E�� ��tH�E�H��H��4������H��Ѕ�u&H�E�� ��t%H�E�H��H��4������H��Ѕ�t
�   �A  H�E�H�PH�E�H�@H��H��H�01������H���H��I��H��w������H���H�U�H�BH�E�H�@H��u
�   ��  H��
      H�H�P�H��
      H��  H��
      H�H��� ��t3H��
      H�H��H��H�
3������H��Ѕ�t
�   �v  H��
      H�H���@H��
      H�H��H���������(W��@�-  H��
      H�H��� ��u�   ��   H��
      H�H�����  H������� ���E�H������H��
      H�H��� ����  �E�H�H������  H������� ���E�H������H��
      H�H��� ���[  �E�H�H������J  H������� ��H��H������F  H������� ���   H)�H��H������"  H������� ���E�H������H��
      H�H�P�H��
      H�H��
      H�� ����  �E�H�H������  H������� ���E�H������H��
      H�H�P�H��
      H�H��
      H�� ���b  �E�H�H��H������N  H��
      H�H�P�H��
      H��6  H��
      H�H��H�E��H�m�H�E؋ ��u�H�E�H��� ����   H���������H��     H�E�H��H�@H�E�H�E�H�P�H������H�BH��
      H�H��D      H�H)�H��H���H*�H�E��@H�E�H�PH��
      H�H�E�H������H��
      H�H��D      H�H)�H��H��H��H����6  H���������H�<I��H��������H��и   �  H�E�H��� ����  H���������H��     H��
      H�H��D      H�H)�H��H���H*�H�E��@H�E�H�PH��
      H�H��
      H�H��
      H�H)�H��H���E�H�E�H��H�@��H��
      H�H��
      H�H)�H��H���E�)ЉE�H��
      H�H�P�H��
      H�H��
      H�H���@�,�H�H��H��H��D      H�H�H��
      H��E�    �_H��
      H��U�Hc�H��H��H�H��
      H�H�PH� H�H�QH��
      H�H�PH��
      H��E��E�;E�|��Z  H���������H�<I��H��!������H��и   �<  H������H�PH������� ���E�H��
      H�H��
      H�H)�H��H���E�)ЉE�H��
      H�H�P�H��
      H�H��
      H�H�� H�@H������H��
      H�H���@�,�H�H��H��H��D      H�H�H��
      H��E�    �_H��
      H��U�Hc�H��H��H�H��
      H�H�PH� H�H�QH��
      H�H�PH��
      H��E��E�;E�|���   �    ��   H������� ���E�H������H������� ���E�H�������UȋẺ։�I��H�� ������H��Ѕ���   �   �   H������� ��H���������H��H�������fI��H�o!������H����RH���������H�<I��H��������H��и   �0��O�����I�����C�����=�����7�����1�����+�����%���H��  [A\A_]���UH��AWSH����H�����I���     L�H��
      H�H��H�E��H�E�H��I��H�t������H���H�m�H��D      H�H9E�sΐ�H��[A_]���UH��AWSH����H�����I��     L�H�}�H�E�H��I��H��������H��Ѕ�t�   �FI��H��������H��Ѕ�tI��H��������H��и   �I��H��������H��и    H��[A_]���UH��AWSH����H�����I��     L�H�}�H�E�H��I��H�������H��Ѕ�t�   �"I��H��������H��Ѕ�t�   ��    H��[A_]���UH��AWATSH��8��H�����I��     L�H�}��u�H�p�������H�L� H�E�H��I��H��m������H���Hc�H��H�H�H��L�H�PH�@H�E�H�UȋE���t
�   �  �E�   �VH��
      H��U�Hc�H��H��H�H��
      H��M�Hcɾ   H)�H��H��H�H�PH� H�H�Q�E��E�;E�~�H��
      H�H�P H��
      H�H��
      H��U�Hc�H��H������H)�H��H��     H��
      H��U�Hc�H��H������H)�H��H�H�E�H�U�H�H�QH��������H�<H�<6������H���H��8[A\A_]���UH��H����H�����I�c�     L؉}��}� ~1�U�Hc�H��
      H�4H��
      H�H)�H��H��H9�~�    �H��
      H��U�Hc�H��H��H�����UH��SH����H�����I�ܢ     L�H�}�H�E� ��t+H�E�H��H�
3������H��Ѕ�tH���������f���	H�E��@H��[]���UH��H����H�����I�n�     L�H�}�H�U����t"H�U�H��H��4������H��Ѕ�t�    �H�E�H�@����UH��AWSH����H�����I��     L�H�}�H�E� ��t"H�E�H��H��4������H��Ѕ�t�    �H�E�H�@H��I��H�P������H���H��[A_]���UH��H����H�����I���     L�H�}�H�E�� ��t�    �H�E�H�@����UH��H����H�����I�M�     L�H�}�H�E�� ��t�    �H�E�H�@����UH��AWSH�� ��H�����I��     L�H�}�H�u�H�E؋ ��t�    �[�E�   H�E�H��H�@2������H���H��I��H��w������H���H�E�H�E�H�@H�U�H��H��I��H��������H���H�� [A_]���UH��AWH��(��H�����I�b�     L�H�}��E�H�U؋��t�    �5�E�   �E��E�H�U�H�RH�M�H��H��I��H��������H���H��(A_]���UH��AWSH�� ��H�����I��     L�H�}�H�E�H��I��H��m������H��ЉE�}� y�    �+H�p�������H�H��E�Hc�H��H�H�H��H�H��H�� [A_]���UH����H�����I�b�     L�H��
      H�H��
      H�H9�w�    �.H��
      H�H�J�H��
      H�H��
      H�]���UH��AWH����H�����I��     L�H��
      H�H��D      H�H)�H��H���  ~'H���������H�<I��H��������H��Ҹ   �H��
      H��    �    H��A_]���UH��AWH����H�����I�K�     L��E�H��
      H�H��D      H�H)�H��H���  ~'H���������H�<I��H��������H��Ҹ   �CH��
      H��   H��
      H�H�JH��
      H�0�E��B�    H��A_]���UH��AWATSH����H�����I���     L�H�}�H��
      H�H��D      H�H)�H��H=�  ~'H���������H�<I��H��������H��и   �nH��
      H��    H�E�H��H�@2������H���H��H��
      L�$I�D$H��
      H�H��I��H��w������H���I�D$�    H��[A\A_]���UH��AWH����H�����I���     L�H�}�H��
      H�H��D      H�H)�H��H���  ~'H���������H�<I��H��������H��Ҹ   �AH��
      H��   H��
      H�H�JH��
      H�0H�E�H�B�    H��A_]���UH��AWH����H�����I�Ǜ     L�H�}�H��
      H�H��D      H�H)�H��H���  ~'H���������H�<I��H��������H��Ҹ   �AH��
      H��   H��
      H�H�JH��
      H�0H�E�H�B�    H��A_]���UH��AWH����H�����I��     L�H�}�H��
      H�H��D      H�H)�H��H���  ~'H���������H�<I��H��������H��Ҹ   �7H��
      H�H�QH��
      H�0H�E�H�PH� H�H�Q�    H��A_]���UH��AWSH�� ��H�����I�F�     L�H�}�H�E�H��I��H��m������H��ЉE�}� y
�   �   H��
      H�H��� ��u�   �iH��
      H�H�P�H��
      H�H��
      H�H�p�������H�H�0�E�Hc�H��H�H�H��H�H�H�QH�FH�V�    H�� [A_]���UH��AWSH��0��H�����I�^�     L�H�}�H�u�H�Eȋ ��t
�   ��   �E�   H�E�H��H�@2������H���H��I��H��w������H���H�E�H�E�H�@H�U�H��H��I��H��������H���H�E�H�}� u�   �dH��
      H�H��� ��u�   �EH��
      H�H�P�H��
      H�H��
      H�H�M�H�PH� H�H�Q�    H��0[A_]���UH��AWSH��0��H�����I�@�     L�H�}��E�H�Eȋ ��t
�   �   �E�   �E��E�H�E�H�@H�U�H��H��I��H��������H���H�E�H�}� u�   �dH��
      H�H��� ��u�   �EH��
      H�H�P�H��
      H�H��
      H�H�M�H�PH� H�H�Q�    H��0[A_]���UH��H����H�����I�J�     L�H�}�H�}� tH�E�� ��u�   ��    ����UH��H����H�����I��     L�H�}�H�}� tH�E�� ��u�   ��    ����UH��H����H�����I���     L�H�}�H�}� tH�E�� ��u�   ��    ����UH��H����H�����I�r�     L�H�}�H�}� tH�E�� ��u�   ��    ����UH��H����H�����I�*�     L�H�}�H�}� tH�E�� ��u�   ��    ����UH��H����H�����I��     L�H�}�H�}� tH�E�� ��u�   ��    ����UH��SH����H�����I���     Lۿ   H��\������H���H�E�H���������H�H�H�E� ��H��H�H� H��H�ob������H��АH��[]���UH��SH����H�����I��     Lۿ   H��\������H���H�E�H�E�H��H��3������H���H��H��d������H��АH��[]���UH��AWSH����H�����I���     L��E�   �-  H�E�H��H��h������H��Ѕ�tEH�E�H��H�]������H����Z�H�8�������H�<I�߸   H�2r������H�����  H�E�H��H�:i������H��Ѕ�tDH�E�H��H��]������H���H��H�<�������H�<I�߸    H�2r������H����n  H�E�H��H��i������H��Ѕ�tDH�E�H��H�c^������H���H��H�@�������H�<I�߸    H�2r������H����  H�E�H��H�j������H��Ѕ�tDH�E�H��H��^������H���H��H�O�������H�<I�߸    H�2r������H����   H�E�H��H��i������H��Ѕ�t.H�E�H��H�]�������H�<I�߸    H�2r������H����gH�E�H��H��h������H��Ѕ�t'H�h�������H�<I�߸    H�2r������H����%H�m�������H�<I�߸    H�2r������H��ҋE�P�U��H��\������H���H�E�H�}� �������H��[A_]���UH��AWATSH��(��H�����I��     L�H�}��E�    �SH��
      H��E�Hc�H��H�H�H��H�H�H�E�H��H��I��H�`E������H��Ѕ�u�E��^  �E�H�����������9E�|�H���������f=�v*H���������H�<I��H��������H��и�����  H��
      H�H�����������H��H�H�H��L�$H�E�H��I��H�P������H���I�$H��
      H�H�����������H��H�H�H��H�H� H��u'H��������H�<I��H��������H��и�����[H��
      H�H����������PH��������f�3��H��H�H�H��H��@   H�������������H��([A\A_]���UH��AWSH��0��H�����I�(�     L�H�}�H�E�H��I��H��H������H��ЉE�E�   ��I��H�4�������H���H�E�H�E��E�   �E�    ��   �E�Hc�H�E�H�� <\��   �E��E�Hc�H�E�H�� ����tt,��tW��nt��rt5�K�E�P�U�Hc�H�E�H�� 
�   �E�P�U�Hc�H�E�H�� 	�|�E�P�U�Hc�H�E�H�� �d�E�P�U�Hc�H�E�H�� \�E�Hc�H�E�H��E�P�U�Hc�H�E�H����&�E�Hc�H�E�H��E�P�U�Hc�H�E�H����E��E��9E�������E�P�U�Hc�H�E�H��  �E�    �gH��      H��U�Hc�H��H�H�H�E�H��H��I��H�`E������H��Ѕ�u%H�E�H��H��I��H���������H��ЋE��   �E�H�����������9E�|�H���������f=� v'H�(�������H�<I��H��������H��и�����SH��      H�H����������PH��������f�3��H��H�H�E�H�H�������������H��0[A_]���UH��AWATSH��(��H�����I�m�     L�H�}��E�    �JH��      H��U�Hc�H��H�H�H�E�H��H��I��H�`E������H��Ѕ�u�E��  �E�H�����������9E�|�H���������f=� v*H�(�������H�<I��H��������H��и�����   H�E�H��I��H��H������H��Ѓ��   ��I��H�4�������H���H�E�H�E�H��      H�H����������PH��������f�3��H��L�$H�U�H�E�H��H��I��H��E������H���I�$H�������������H��([A\A_]���UH��AWH����H�����I��     L�H�}�H�U���uH�E�H�@H��� �7H�U���u,H�U�H�R���uH�U�H�RH��I��H�������H��ҐH��A_]���UH��SH����H�����I�^�     L��E�    �?H��
      H��E�Hc�H��H�H�H��H�H��H��H�t������H��ЃE�H�����������9E�|���H��[]���UH��AWSH����H�����I�Њ     L�I��H�XY������H���H��t������H����E�    �E�E���   H�       H��U�Hc�H��H�H� H��� <ujH�       H��U�Hc�H��H�H�       H�4�E�P�U�H�H��H�H�H�H�       H��U�Hc�H��H�H� H���  �7H�       H��U�Hc�H��H�H� H��H��I��H���������H��ЃE�H��U      ���9E������E��H��U      f��E�    �E��E���   H�      H��U�Hc�H��H�H� � <ufH�      H��U�Hc�H��H�H�      H�4�E��P�U�H�H��H�H�H�H�      H��U�Hc�H��H�H� �  �3H�      H��U�Hc�H��H�H� H��I��H�������H��ЃE�H��U      ���9E��$����E���H��U      f��H��[A_]���UH��AWSH����H�����I�o�     L�H�}�H�}� u
�    �   H��U      �f=�vKH�!u������H���H��U      �f=�v'H�L�������H�<I��H��������H��и    �CH�       H�H��U      ��PH��U      f�3��H��H�H�E�H�H�E�H��[A_]���UH��AWSH����H�����I���     L�H�}�H�}� u
�    �   H��U      �f=�vKH�!u������H���H��U      �f=�v'H�b�������H�<I��H��������H��и    �CH�      H�H��U      ��PH��U      f�3��H��H�H�E�H�H�E�H��[A_]���UH��AWATSH����H�����I���     L�H�}�H��     ���~*H�y�������H�<I��H��������H��и   �   H��     D�$A�D$H��     �H�E�H��I��H�P������H���H�8�     Ic�H�H��H�8�     Ic�H�H��H��u'H��������H�<I��H��������H��и   ��    H��[A\A_]���UH����H�����I���     L�H��     ���H�8�     Hc�H�H��]���UH��AWSH�� ��H�����I�U�     Lۿ   I��H��\������H���H�E�H�}� u%H���������H�<I��H��������H����~  �   I��H��\������H���H��t%H���������H�<I��H��������H����=  H�E�� ��u�E�    �m  H�E�� ��t%H���������H�<I��H��������H�����  �E�    �OH�E�H�HH��
      H�4�E�Hc�H��H�H�H��H�H� H��H��I��H�`E������H��Ѕ�t�E�H�����������9E�|���H�����������9E�u%H��������H�<I��H��������H����J  �E���E�H�������������9E�},H��
      H��E�Hc�H��H�H�H��Hȋ@��t�H�������������9E�u)I��H�a������H���I��H�a������H����   �E�   H��
      H��E�Hc�H��H�H�H��H�H� H��I��H�@2������H���H��H��w������H���H�E�H�E�H��I��H��d������H��Ѕ�uAH��
      H��E�Hc�H��H�H�H��H�H��H��I��H��d������H��Ѕ���H�� [A_]���UH��AWSH����H�����I�`�     Lۉ��E�H��      H�H�ص      H�H)�H��H=�  ~1H�8�������H�<I��H��������H���H� �      �   H��      H�H�PH��      H��U��H��[A_]���UH��AWSH����H�����I���     Lۉ�f�E�H��      H�H�ص      H�H)�H��H=�  v1H�8�������H�<I��H��������H���H� �      �   H��      H��U�f�H��      H�H�PH��      H��H��[A_]���UH��AWSH����H�����I��     L��E�H��      H�H�ص      H�H)�H��H=�  v1H�8�������H�<I��H��������H���H� �      �   H��      H��E�� H��      H�H�PH��      H��H��[A_]���UH��AWS��H�����I��     L�H��      ���H��      �Ѓ�^H��      ��PH��      ��1H�M�������H�<I��H��������H���H� �      �   �[A_]���UH��AWS��H�����I��     L�H��      ���H��      �Ѓ�^ H��      ��PH��      ��1H�`�������H�<I��H��������H���H� �      �   �[A_]���UH��AWS��H�����I��~     L�H���      �<w H���      ��PH���      ��1H���������H�<I��H��������H���H� �      �   �[A_]���UH��SH����H�����I�S~     Lۉ}�}�v�E�   ��    H��}������H���H��      H�H�PH�      H�H)�H�ЋM�H�H��H��H��u���H��[]���UH��SH��(��H�����I��}     L��E��E��,��E��*E�.E���   .E���   �}� �E������H��}������H�����   �}��   2�   H��}������H��ЋE�����H��}������H����   �   H���������H��п   H��}������H��ЋE�����H�H~������H����A�   H���������H��п   H��}������H��ЋE�fn�H�������H���H��������H��АH��([]���UH��H����H�����I�||     L؉�f�U�H��      ��҃��U��&H��      �U�Hc�H��Qf9U�u�E���m��}� yԸ��������UH��SH����H�����I�|     L�H�}�H�}� ~[�   H���������H��п   H��}������H���H�E������H�H~������H���H��������H����   H�}� yiH�U�H�}�	H�E��	����H��}������H����.�   H��}������H���H�E�����H��}������H���H��������H����2�   H��}������H���H��      ��P�H��      ��H��[]���UH��SH����H�����I��z     Lۉ}�'   H��}������H��ЋE��H��      ������H��}������H��АH��[]���UH��SH��(��H�����I�az     Lۉ}�H���      �E�H�H�H��H��~]�   H���������H��п#   H��}������H���H���      �E�H�H�H������H�H~������H����1  H���      �E�H�H�H��H��ysH���      �E�H�H�H���ЉE��}�	 �E�������H��}������H�����   �"   H��}������H��ЋE�����H��}������H����   �E�    �E܃��E��#H���      �E�H�H�H��H��u�E��E�H���      ���9E�|ǋE� �E�ЉE�}� u�$   H��}������H����-�%   H��}������H��ЋE�����H��}������H��АH��([]���UH��AWAUATSH����H�����I��x     L�H�}�I��H�Vz������H���I��H���������H�D�(I��H�l%������H���H��H�E�M��E��H��H��H���������H�4H�X�      H�<I�߸    I�in������I�A��H�X�      H�<I��H��������H���H� �      �   �H��[A\A]A_]���UH����H�����I��w     Lظ   ]���UH��AWSH����H�����I�rw     L�H�      H�H�E�H� �      �    �    H�b�������H��҅�uH� �      ���u�   �^H�      H�H�PH�      H�� <H�E�H��I��H�<6������H��Ѕ�t�   �H�      H�E�H��    H��[A_]���UH��AWAVAUATSH��H��H�����I��v     L��E̖   �E�����I��H��������H���H�(�      H��E�����I��H��������H���H�0�      H�H�(�      H�H��tH�0�      H�H��u(H���������H�<H�k�������H��и   �?!  H�(�      H�H�P�H�8�      H�H�0�      H�H�P�H�@�      H�H�H�      �    H�L�      �    H���     �    H���     �    H���     ������H�8�      H�H�E�H�@�      H�H�E�H�H�      D�4H�E�H�u�H�u�H�0�      H��U�H��H�H9��~  H�0�      H�H)�H��H���E�H�(�      H�H�u�H)�H��H���E�H�(�      H�I)�L��H���E��E̖   �E̍�    H�(�      H���H��I��H�υ������H���H�(�      H��E̍�    H�0�      H���H��I��H�υ������H���H�0�      H�H�(�      H�H��tH�0�      H�H��u(H���������H�<H�k�������H��и   �%  H�0�      H��U�Hc�H��H�H�E�H�(�      H��U�Hc�H��H�H�E�H�(�      H��U�Hc�H��L�$H�E�D�0H�E�H�u�H�u�H���     H�H�H�ؽ������Ic�H�D�,�A������  H���     ���yFI�߸    H��%������H���H���     �H���     ���yH���     �    H���     �A�E����   A��=  ��   H�ظ������Ic�H�D�,�H���������Ic�Hڋ�H���     �9�umH���     �����H���     H���     H�H�E��H���     �������H���     ��P�H���     �����������H���������Ic�H�D�,�A�����   H���     ���yFI�߸    H��%������H���H���     �H���     ���yH���     �    H���������L�,�I��A�E ���u�I�E� A9�u�I��A�E ��xA�U H���     �9�u�E�mE��yPH�0�      H�H��I��H���������H���H�(�      H�H��I��H���������H��и    �J  E����  H���     ����9  ����  ��t����  ������  �H���������H�<H�k�������H��АH���     �   �|H�E�� H�ؽ������H�Hڋ�D��   E��xNA��=  EH�ظ������Ic�Hڋ�H���������H�Hڋ�=   uH�ظ������Ic�H�D�4������H�m�H�m�H�0�      H�H9E��l���H�0�      H�H��I��H���������H���H�(�      H�H��I��H���������H��и   ��  H���     ���uPH�0�      H�H��I��H���������H���H�(�      H�H��I��H���������H��и   �  H���     ����������H�L�      D�,H�u�I��H�8�������Ic�H�D�4�D��������   A��Ic�H��H��H�H�u�H���     H�FH�H�x�������Ic�H�D�,�H���������Ic�Hڋ�Ic�H��H��HE�H�M�H�M���D�pA��=  4H�ظ������Ic�H�D�4�H���������Ic�Hڋ�D����9��%���H���������Ic�Hڋ�H�ظ������H�H�D�4������A��Ic�H��H��HE�H�u�H�u�H���     H�FH�H�x�������Ic�H�D�,�H���������Ic�Hڋ�Ic�H��H��HE�H�M�H�M���D�pA��=  0H�ظ������Ic�H�D�4�H���������Ic�Hڋ�D����9�t&H���������Ic�Hڋ�H�ظ������H�H�D�4�H�H�      D�4H�@�      H�M�H�H�8�      H�u�H�4H�L�      ���h�������H��    H��R H�H��R H�>��H�      H�H�ص      H�H�ص      H�H��      H�H��      � ��  H��      H�H�      H���  H�      H�H�ص      H�H�ص      H�H��      H�H��      � �|  H�x�������H�� ��td�   H���������H��п=   H��}������H���I�D$�� ����H�H~������H���I�D$�� ����H�H~������H��п    H�#�������H�����  H�x�������H�� ��t�?   H��}������H��п;   H��}������H���H��      �����H��}������H���H�p�������H�H�I�D$�� ��H��H�H�H��H��@   H��      H�H�      H�H)�H�Љ�H�p�������H�H�I�D$�� ��H��H�H�H��L�,�   I��H�4�������H���I�EH��      H�H�      H�H)�H�Љ�H�      H�H�p�������H�H�0I�D$�� ��H��H�H�H��H�H�@��H��H��I��H��B������H����i  H��      �    H�x�������H�� ���  �   H���������H��п>   H��}������H���H���������H�� ����H�H~������H�����  I�D$�H� H��H�E�H��      H�H9E�u4H��      H�H�P�H��      H�H��      H�H�E��/I�D$�H� � 5H��      H�H+E�H��I�D$�H� H��f�I�D$�H� � 7I�D$�H� H�PH�E�H)�H��I�D$�H� H��f��0  H��      H�H���     H��  I�D$�H� � 7H��      H�I�D$�H� H��H)�I�D$�H� H��f�I�D$�H� � 6H��      H�I�D$�H� H)�I�D$�H� H��f��  H��      H�H���     H��  I�$� 8H��      H�I�D$�H� H)�I�$H��f��O  A�$��t/H���      ���H��      �I�D$�� �)���9�t/I�D$�� � H���      ���Љ�H�#�������H���H���      ������E���E���H���������H��Ѓm��}� y�I�D$�� ��'I�D$�� ���p  H���      H�H���Y  �    H�#�������H����?  �    H�#�������H����J  I�D$�H� H��H�E�H��      H�H9E�u4H��      H�H�P�H��      H�H��      H�H�E��/I�D$�H� � 5H��      H�H+E�H��I�D$�H� H��f�I�D$�H� � 7I�D$�H� H�PH�E�H)�H��I�D$�H� H��f��  H��      ���H���     ��k  H��      �    �U  H��      ���I�D$� 9��  I�D$� ��H��      ��    H�#�������H�����  H�x�������H�� ����  �   H���������H��п>   H��}������H���H���������H�� ����H�H~������H����  H�x�������H�� ��t�?   H��}������H��п;   H��}������H���H��      �����H��}������H����3  �   H���������H���H��      H�H���     H��    H��}������H��п    H�H~������H�����  A�$����  H��      �����H�#�������H���H��������H����}  I�D$�� H���     ��w  �)   H��}������H���H���     �   H��      ��P�H��      ��/  �*   H��}������H���H���     �   H��      ��P�H��      ���  �+   H��}������H��п2   H��}������H���H���     �   H��      ��P�H��      ��  �)   H��}������H��п2   H��}������H���H���     �   H��      ��P�H��      ��-  �+   H��}������H���H���     �   H��      ��P�H��      ���  �*   H��}������H��п2   H��}������H���H���     �   H��      ��P�H��      ��  �,   H��}������H���H���     �   H��      ��P�H��      ��@  �-   H��}������H���H���     �   H��      ��P�H��      ���  �.   H��}������H���H���     �   H��      ��P�H��      ��  �/   H��}������H���H���     �   H��      ��P�H��      ��h  �0   H��}������H���H���     �   H��      ��P�H��      ��   H���     �   �
  �1   H��}������H���H���     �   ��  �   H��}������H���H��      H�H���     H��    H��}������H���H��������H��п(   H��}������H����o  A�$I�D$�H� �I�D$�H� H��yH���     �   �1  I�D$�H� H��H��H��������H��п   H��}������H���H��������H��п   H��}������H���H��������H��п:   H��}������H���H��      ��P�H��      �H���     �    H�x�������H�� ���m
  �   H���������H��п>   H��}������H���H���������H�� ����H�H~������H����
  �(   H��}������H���H���     �   ��	  I�$H��H��������H���H���     �   ��	  A�$fn�H�+�������H���H���     �   �	  �   H���������H��п   H��}������H���A�$����H�H~������H���H���     �   H��������H����6	  �   H��}������H���H���     �   H��������H�����  H���     �    H�x�������H�� ����  �   H���������H��п>   H��}������H���H���������H�� ����H�H~������H����w  �2   H��}������H���H���     �   �S  �9   H��}������H���H��      ��P�H��      ��  I�D$�H� � 4H��      H�I�D$�H� H��H)�I�D$�H� H��f�H���     �   ��  �9   H��}������H���H��      ��P�H��      ��  I�D$�H� � 3H��      H�I�D$�H� H��H)�I�D$�H� H��f�H���     �   �K  �   H��}������H���H��������H����!  �   H��}������H���H��      �H���     �H��������H�����  �:   H��}������H���I�D$� �P�H��      ��  I�$H��H��������H����  H���     �   �z  A�$H���     ��d  A�$H���     ��N  I�D$�� ���>  H��      �����H�#�������H���H��������H����  A�$H���     ���  H��      ���A�$H��      H�H�f�AH�u�������H����  H��      ���A�$H��      H�H�f�AH�u�������H����v  H���     H������_  A�$��H���     H��D  I�D$�� H���     ��+  I�D$�� H���     ��  H���     �    ��  A�$H���     ���  H���     �   ��  I�D$�� �PH���     ��  �   H���������H��п   H��}������H���H�p�������H�H�A�$��H��H�H�H��H�H� H��I��H��r������H�������H�H~������H���H��������H����  �&   H��}������H���H��      ��P�H��      ���  H���     �    ��  A�$H���     ��  H�P��������H�+�������H����  H���     �   �  I�D$�� ���*�H�+�������H����_  I�D$� �PH���     ��C  �&   H��}������H���H��      ��P�H��      ��  H���      � H���      ���I�$H���      H�H�H��H��������H���I�$H������H���     ��  H���      ���I�$H���      H�H�H��H��������H���I�$H��uI�D$�� ���I�D$�� H���     ��A  A�$����H�x�������H��ЉE��}��u A�$����H�H���     H���  �E���H�H���     H���  I�$H��H��������H�����  H���     H�    �  I�$H��H��������H����  �   H���������H��п   H��}������H���H�p�������H�H�A�$��H��H�H�H��H�H� H��I��H��r������H�������H�H~������H���H��������H���H���     H�    ��   I�D$�H��      ����H��      Hc�H�3f�AH�u�������H����   I�D$�H��      ����H��      Hc�H�3f�AH�u�������H����k�   H��}������H����TH��      �    �AA�$H�x�������H���+�������{�����u�����o�����i�����c�����]�����W���H��H[A\A]A^A_]���UH��AWS��H�����I�sT     Lۿ   I��H��\������H���H��I��H��d������H��о   H�X�������H�<I��H��Z������H��А[A_]���UH��AWSH����H�����I��S     Lۿ   I��H��\������H���H�E�H�E�H��I��H�:i������H��Ѕ�t3H�E�H��I��H��]������H��о    H��I��H��Z������H��АH��[A_]���UH��AWSH����H�����I�YS     Lۿ   I��H��\������H���H�E�H�E�H��I��H�:i������H��Ѕ�t.H�E�H��I��H��]������H���H��I��H�rZ������H��АH��[A_]���UH��AWSH�� ��H�����I��R     Lۉ}�H�u�H���������H�H�H�X�������H�H�H�8�������H�H�H���������H�H�H���������H�H�H���������H�H�H�8�������H�H�H���������H�H��}�%H�`�������H�<I��H��q������H����\  H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���I��H���������H���I��H���������H���I��H���������H���H�E�H��H� H��I��H��Y������H����E�   �5�E�H�H��    H�E�H�H� �    H��I��H��Z������H��ЃE��E�;E�|�H�� [A_]���UH��AWSH����H�����I�|P     Lۿ   I��H��\������H���H�E�H�}� ��   H�       H�H���������H�H� H9�tBH�       H�H��I��H��S������H���H���������H�H� H�       H�H����������I��H��a������H����E  H�E�H��I��H�:i������H��Ѕ�uEH���������H�<I��H��������H���H���������f��I��H��a������H�����   H�E�H��I��H��]������H���H���������H�4H��I��H�VS������H���H�E�H�}� u"H���������f��I��H��a������H����zH�       H�H���������H�H� H9�t#H�       H�H��I��H��S������H���H�       H�E�H�H����������I��H��a������H��АH��[A_]���UH��AWSH����H�����I�TN     Lۿ   I��H��\������H���H�E�H�}� ��   H�      H�H�8�������H�H� H9�tBH�      H�H��I��H��S������H���H�8�������H�H� H�      H�H����������I��H��a������H����E  H�E�H��I��H�:i������H��Ѕ�uEH���������H�<I��H��������H���H���������f��I��H��a������H�����   H�E�H��I��H��]������H���H���������H�4H��I��H�VS������H���H�E�H�}� u"H���������f��I��H��a������H����zH�      H�H�8�������H�H� H9�t#H�      H�H��I��H��S������H���H�      H�E�H�H����������I��H��a������H��АH��[A_]���UH��AWSH��  ��H�����I�)L     Lۿ   I��H��\������H���H�E�H�}� �  �H�       H�H��I��H��U������H��ЉEЋE���H���������H�H������ ��u��}�"u]H�       H�H������H���������H�4H��I�߸    H�}������H��у��N  I��H�a������H����  �}�'u]H�       H�H������H��������H�4H��I�߸    H�}������H��у���   I��H�a������H����O  H�       H��E�H�։�I��H��~������H���H�       H�H������H�	�������H�4H��I�߸    H�}������H��у�tI��H�a������H�����  H�U�H������H��H��I��H�̓������H���fH~�H�E�H�E�� ��u�ZE�I��H��a������H����{  H������H��I��H�ob������H����Z  H�E�H��I��H��]������H���H�E��E�    �H�E�H�E�� ��H���������H�H������ ��u�H�E�H�PH�U�� �E��(�U��������H�E�H�PH�U�� ����0ȉE�H�E�� ��H���������H�H��������u��}� �`  �U�H��P���H��������H�4H��I�߸    H�in������H���H�       H�H������H��P���H��H��I�߸    H�}������H����E׉�I��H�
R������H��Ѓ�g
��e}a�   ��i��   H�U�H������H��������H�4H��I�߸    H�'s������H���H�E��H*�I��H��a������H����  H�U�H������H��������H�4H��I�߸    H�'s������H��ыE�fn�I��H��a������H����Z  H������H��I��H�ob������H����9  �E׉�I��H�
R������H��Ѓ�g
��e}h�   ��i��   H�       H�H�U�H��������H�4H��I�߸    H�}������H���H�E��H*�I��H��a������H����   H�       H�H�U�H��������H�4H��I�߸    H�}������H��ыE�fn�I��H��a������H����ZH�       H�H������H�	�������H�4H��I�߸    H�}������H���H������H��I��H�ob������H��АH�Ġ  [A_]���UH��AWATSH��H��H�����I�nF     L�H�}�H�u�H�W�      H�H�E��E�r�E�    �E�    �H�E�H�E�� ��H���������H�H������ ��u�H�E�H�PH�U�� �E�H�E�� <<tH�E�� <|tH�E�� <>u<H�E�H�PH�U�� �E��(�UЉ�������H�E�H�PH�U�� ����0ȉE�H�E�� ��H���������H�H��������u�H�E��(�Ủ�������H�E�H�PH�U�� ����0ȉE�H�E�� ��H���������H�H��������u�H��������H�4H�X�      H�<I�߸    H�in������H��Ҁ}�<t�}�|uM�    H�X�      H�<I��H��D������H���H��������H�4H��I�߸    H�in������H��҃}� tU�    H�X�      H�<I��H��D������H���H���EЉ�H��������H�4H��I�߸    H�in������H��у}� tU�    H�X�      H�<I��H��D������H���H���Ẻ�H�!�������H�4H��I�߸    H�in������H���D�eþ    H�X�      H�<I��H��D������H���D��H�%�������H�4H��I�߸    H�in������H����EÉ�I��H�
R������H��Ѓ�s��   ��s�  ��g
��e}a��   ��i��   �E�iH�E�H��I��H�]������H����H,�H�E�H�X�      H�4H��I�߸    H�in������H����   �E�fH�E�H��I��H�]������H����Z�H�E�H�X�      H�4H��I�߸   H�in������H����a�E�sH�E�H��I��H��]������H���H��H�E�H�X�      H�4H��I�߸    H�in������H����H�(�������H��  H�E�H��I��H��H������H��ЉE��}� tB�E�;E�~:�E�    ��E�Hc�H�E�H�� *�E��E�;E�|�E�Hc�H�E�H��  �   �}� ��   �}�|��   �E����E���m��E�Hc�H�E�H�� ��H���������H�H������ ��uˋE�+Eĉ������H�H��HE��E�    ��EčP�U�Hc�H�E�H��  �E�Hc�H�E�H�� ��t֋E�Hc�H�E�H��  H�E�H��H[A\A_]���UH��AWSH�� ��H�����I� A     Lۿ   I��H��\������H���H�E�   I��H��\������H���H�E�H�}� u\H�      H�H�)�������H�4H��I�߸    H��c������H���H����������I��H��a������H�����  H�}� �
  �E�    H�E�H��I��H��h������H��Ѕ�tXH�E�H��I��H�]������H����Z�H�      H�H�+�������H�4H��I�߸   H��c������H��҉E��rH�E�H��I��H�:i������H��Ѕ�tUH�E�H��I��H��]������H���H��H�      H�H�	�������H�4H��I�߸    H��c������H��щE��*E�I��H��a������H�����   H�E�H��I��H�:i������H��Ѕ�uEH�0�������H�<I��H��������H���H���������f��I��H��a������H����   H�E�H��I��H��]������H���H��H�E�H��H��H���������H���H��H�      H�H�	�������H�4H��I�߸    H��c������H����*�I��H��a������H���H�� [A_]���UH��AWSH����H�����I�;>     Lۿ   I��H��\������H���H�E�H�}� tH�E�H��I��H�:i������H��Ѕ�uBH�X�������H�<I��H��������H���H���������f��I��H��a������H����OH�E�H��I��H��]������H���H��I��H�p�������H���H����������I��H��a������H��АH��[A_]���UH��AWSH����H�����I�:=     Lۿ   I��H��\������H���H�E�H�}� tH�E�H��I��H�:i������H��Ѕ�uBH�X�������H�<I��H��������H���H���������f��I��H��a������H����uH�E�H��I��H��]������H���H��I��H��X������H��Ѕ�u#H����������I��H��a������H����!H���������f��I��H��a������H��АH��[A_]���UH��AWS��H�����I�<     L�H�u�������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H�ų������H�<I��H�fc������H���H���������H�<I��H��e������H���H��������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H��А[A_]���UH��AWSH����H�����I�j:     Lۿ   I��H��\������H���H�E�H�}� u%H���������H�<I��H��������H����   H�E�H��I��H��h������H��Ѕ�u"H���������H�<I��H��������H����kH�E�H��I��H�]������H����Z��E�H��������f��f/E�v�E�H��������f(fW��E��ZE�I��H��a������H���H��[A_]���UH��AWSH����H�����I�I9     Lۿ   I��H��\������H���H�E�H�}� u%H��������H�<I��H��������H����   H�E�H��I��H��h������H��Ѕ�u"H�0�������H�<I��H��������H����SH�E�H��I��H�]������H����Z��E�H�E�fHn�I��H��������H����Z�I��H��a������H���H��[A_]���UH��AWSH����H�����I�@8     Lۿ   I��H��\������H���H�E�H�}� u%H�X�������H�<I��H��������H����   H�E�H��I��H��h������H��Ѕ�u"H���������H�<I��H��������H����SH�E�H��I��H�]������H����Z��E�H�E�fHn�I��H���������H����Z�I��H��a������H���H��[A_]���UH��AWSH����H�����I�77     Lۿ   I��H��\������H���H�E�H�}� u%H���������H�<I��H��������H����   H�E�H��I��H��h������H��Ѕ�u"H���������H�<I��H��������H����SH�E�H��I��H�]������H����Z��E�H�E�fHn�I��H�R�������H����Z�I��H��a������H���H��[A_]���UH��AWSH����H�����I�.6     Lۿ   I��H��\������H���H�E�H�}� u%H���������H�<I��H��������H����   H�E�H��I��H��h������H��Ѕ�u"H� �������H�<I��H��������H����SH�E�H��I��H�]������H����Z��E�H�E�fHn�I��H�ա������H����Z�I��H��a������H���H��[A_]���UH��AWSH����H�����I�%5     Lۿ   I��H��\������H���H�E�H�}� u%H�H�������H�<I��H��������H����   H�E�H��I��H��h������H��Ѕ�u"H�p�������H�<I��H��������H����SH�E�H��I��H�]������H����Z��E�H�E�fHn�I��H���������H����Z�I��H��a������H���H��[A_]���UH��AWSH����H�����I�4     Lۿ   I��H��\������H���H�E�H�}� u%H���������H�<I��H��������H����   H�E�H��I��H��h������H��Ѕ�u"H���������H�<I��H��������H����SH�E�H��I��H�]������H����Z��E�H�E�fHn�I��H�c�������H����Z�I��H��a������H���H��[A_]���UH��AWSH����H�����I�3     Lۿ   I��H��\������H���H�E�H�}� u%H���������H�<I��H��������H����   H�E�H��I��H��h������H��Ѕ�u"H��������H�<I��H��������H����SH�E�H��I��H�]������H����Z��E�H�E�fHn�I��H���������H����Z�I��H��a������H���H��[A_]���UH��AWSH����H�����I�
2     Lۿ   I��H��\������H���H�E�H�}� u%H�8�������H�<I��H��������H����   H�E�H��I��H��h������H��Ѕ�u"H�`�������H�<I��H��������H����SH�E�H��I��H�]������H����Z��E�H�E�fHn�I��H�Ģ������H����Z�I��H��a������H���H��[A_]���UH��AWSH�� ��H�����I�1     Lۿ   I��H��\������H���H�E�   I��H��\������H���H�E�H�E�H��I��H��h������H��Ѕ�tH�E�H��I��H��h������H��Ѕ�u"H���������H�<I��H��������H����_H�E�H��I��H�]������H����,��E�H�E�H��I��H�]������H����,��E؋Eܙ�}؉��*�I��H��a������H���H�� [A_]���UH��AWSH����H�����I��/     Lۿ   I��H��\������H���H�E�H�}� u%H���������H�<I��H��������H����   H�E�H��I��H��h������H��Ѕ�u"H���������H�<I��H��������H����SH�E�H��I��H�]������H����Z��E�H�E�fHn�I��H�(�������H����Z�I��H��a������H���H��[A_]���UH��AWSH�� ��H�����I��.     Lۿ   I��H��\������H���H�E�   I��H��\������H���H�E�H�E�H��I��H��h������H��Ѕ�tH�E�H��I��H��h������H��Ѕ�u"H� �������H�<I��H��������H����~H�E�H��I��H�]������H����Z��E�H�E�H��I��H�]������H����Z��E��E�H�E�f(�fHn�I��H���������H����Z�I��H��a������H���H�� [A_]���UH��AWSH�� ��H�����I��-     L��E�   �E�P�U��I��H��\������H���H�E�H�}� u%H�(�������H�<I��H��������H����"  H�E�H��I��H��h������H��Ѕ�u%H�P�������H�<I��H��������H�����   H�E�H��I��H�]������H����Z��E��yH�E�H��I��H��h������H��Ѕ�u"H�P�������H�<I��H��������H����}H�E�H��I��H�]������H����Z��E��E�f/E�w�
�E��E��E�P�U��I��H��\������H���H�E�H�}� �[����ZE�I��H��a������H���H�� [A_]���UH��AWSH�� ��H�����I��+     L��E�   �E�P�U��I��H��\������H���H�E�H�}� u%H�x�������H�<I��H��������H����"  H�E�H��I��H��h������H��Ѕ�u%H���������H�<I��H��������H�����   H�E�H��I��H�]������H����Z��E��yH�E�H��I��H��h������H��Ѕ�u"H���������H�<I��H��������H����}H�E�H��I��H�]������H����Z��E��E�f/E�w�
�E��E��E�P�U��I��H��\������H���H�E�H�}� �[����ZE�I��H��a������H���H�� [A_]���UH��AWS��H�����I�O*     L�H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H��������H�<I��H�fc������H���H���������H�<I��H��e������H���H��������H�<I��H�fc������H���H���������H�<I��H��e������H���H�Z�������H�<I��H�fc������H���H���������H�<I��H��e������H���H� �������H�<I��H�fc������H���H��������H�<I��H��e������H��А[A_]���UH��AWSH��0��H�����I��&     Lۿ   I��H��\������H���H�E�   I��H��\������H���H�E�H�E�H��I��H�:i������H��Ѕ�tH�E�H��I��H�:i������H��Ѕ�u"H�(�������H�<I��H��������H����{H�E�H��I��H��]������H���H�E�H�E�H��I��H��]������H���H�E�H�U�H�E�H��H��I��H�jO������H���H+E؃��E��*E�I��H��a������H���H��0[A_]���UH��AWSH����H�����I�e%     Lۿ   I��H��\������H���H�E�H�E�H��I��H�:i������H��Ѕ�u"H�X�������H�<I��H��������H����cH�E�H��I��H��]������H���H��I��H��H������H��Љ�H��x�H*��H��H���H	��H*��X�I��H��a������H���H��[A_]���UH��AWSH��0��H�����I�x$     Lۿ   I��H��\������H���H�E�   I��H��\������H���H�E�   I��H��\������H���H�E�H�E�H��I��H�:i������H��Ѕ�t:H�E�H��I��H��h������H��Ѕ�tH�E�H��I��H��h������H��Ѕ�u%H���������H�<I��H��������H����  H�E�H��I��H��]������H���H��I��H�P������H���H�E�H�E�H��I��H�]������H����,��E�H�E�H��I��H�]������H����,��EȋE�;E�|&�}� ~ H�E�H��I��H��H������H��ЋU�9�s"H���������H�<I��H�ob������H����5�E�Hc�H�E�H��  �E�H�H�P�H�E�H�H��I��H�ob������H���H�E�H��I��H���������H���H��0[A_]���UH��AWSH�� ��H�����I�k"     Lۿ   I��H��\������H���H�E�H�E�H��I��H�:i������H��Ѕ�u%H���������H�<I��H��������H����   H�E�H��I��H��]������H���H��I��H�P������H���H�E�H�E�H�E��+H�E�� ����I��H�
R������H��Љ�H�E�H�E�H�E�� ��u�H�E�H��I��H�ob������H���H�E�H��I��H���������H���H�� [A_]���UH��AWSH�� ��H�����I�:!     Lۿ   I��H��\������H���H�E�H�E�H��I��H�:i������H��Ѕ�u%H���������H�<I��H��������H����   H�E�H��I��H��]������H���H��I��H�P������H���H�E�H�E�H�E��+H�E�� ����I��H�_R������H��Љ�H�E�H�E�H�E�� ��u�H�E�H��I��H�ob������H���H�E�H��I��H���������H���H�� [A_]���UH��AWS��H�����I�      L�H�O�������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H�y�������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H���������H�<I��H��e������H���H���������H�<I��H�fc������H���H��������H�<I��H��e������H��А[A_]���UH��AWSH����H�����I��     Lۉ}�H�u�H�E�� ��H�E��@9�sH�E��P#H�E��@9�r"H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@��u)H�8�������H�H��E�H�։�H�Q�������H���H�E�H�PH�E��@#��H�H�E�H�PH�E�H�@�U�H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  H�E��@��u0H���������H�H� H��t�E�����I��H�5������H��ЋE�H��[A_]���UH��H����H�����I�I     L�H�}��E�    H�E�@��u]H�E�@'�PH�E�P'��H�E�P#H�E�@'9�r�H�E�H�PH�E�@'��H��H�H�E�H�PH�E�H�@� ���E��   H�E�@��tH�E�@��uiH�E�@#��u������ZH�E�P'H�E�@#9�r������AH�E�H�PH�E�@'��H�H�E�H�PH�E�H�@� ���E�H�E�@'�PH�E�P'�E�����UH��H����H�����I�+     L�H���������H�H� H�E��E�    H�E��@��uWH�E��P#H�E��@'9�w�    �AH�E�H�PH�E��@'��H�H�E�H�PH�E�H�@� ���E�H�E��@'�PH�E��P'�E�����UH��H����H�����I��     L�H���������H�H� H�E��E�    H�E��@��uXH�E��@'�PH�E��P'��H�E��P#H�E��@'9�r�H�E�H�PH�E��@'��H��H�H�E�H�PH�E�H�@� ���E��E�����UH��AWH��(��H�����I��     L�H�}�H�u�H�U����u�    �(H�M�H�U�H��H��I��H���������H���H�E�H�E�H��(A_]���UH��AWSH�� ��H�����I�g     L�H�}�H�}� u
������   H�}� tH�E؋@����tH�E��@"<t������zH�E؋@%�   ��u�    �cH�E؋@#H�U؋J�    ��E�H�E؋@��@��u�U�H�E؉�H��I��H�C������H���H�E�H��I��H�5������H��ЉE�E�H�� [A_]���UH��AWSH����H�����I��     L�H�}�H�}� u������0H�E�H��H���������H���H�E�H��I��H�o������H���H��[A_]���UH��AWSH�� ��H�����I�     Lۉ}�H�u�H�}� u
�������  H�EЋ@��u
�    �  H�EЋ@��tH�EЋ@��tH�EЋ@��u!H�UЋE�H�։�H�Q�������H����y  H�EЋ@����unH�EЋP#H�EЋ�+  9�wYH�EЋ�+  ��tKH�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��E�U�H�EЉ�H��I��H�o������H����H�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U܈H�E�� ��H�EЋ@��9�r3H�EЋ@����H�EЉPH�E�f�   H�E�H��H���������H���H�EЋ@#�PH�EЉP#H�EЋP#H�EЋ�+  9�vH�EЋ�+  �PH�EЉ�+  H�EЋ@���H�EЉP�    H�� [A_]���UH��AWH��(��H�����I��     L�H�}�H�}� u
������  H�E؋@��u
�    �v  H�E؋@��tH�E؋@��tH�E؋@��u"H�E�H��H���������H��ЉE�E��0  H�E؋P#H�E؋�+  9�r
������  H�E؋@����ulH�E؋P#H�E؋�+  9�wWH�E؋�+  ��tIH�E؋@����H�E؉PH�E؋@#H�U؋r�    ���E�U�H�E؉�H��I��H�o������H���H�E؋@#H�U؋J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@� ���E�H�E�� ��H�E؋@��9�rH�E؋@����H�E؉PH�E�f�   H�E؋@#�PH�E؉P#�E�H��(A_]���UH��SH��H��H�����I�%     L�H�}ȉuĉU�H�M�H�}� u�    �y�E�    H�E�H�E��E�    �FH�E�H��H���������H��ЉE؃}��u�E�    �u��4H�E�H�PH�U��U؈�E��E��E��E��E�9�w��E�    �u�H��H[]���UH��SH��H��H�����I�d     L�H�}ȉuĉU�H�M�H�}� u�    �l�E�    H�E�H�E��E�    �9H�E�H�PH�U�� ���E�H�U��E�H�։�H���������H��ЃE��E��E��E��E�9�w��E�    �u�H��H[]���UH��H����H�����I��     L�H�}�H�u��U�}�tZ�}�|�}� t�}�t�nH�E���H�E��P#H�E���H�E��P'�RH�E��@#H�U��H�E��P#H�E��@'H�U��H�E��P'�(H�E���+  H�U�)Љ�H�E��P#H�E��P#H�E��P'�H�E��@#H�U��J�    ��Љ�H�E�f��    ����UH��H����H�����I��     L�H�}�H�}� u�    �	H�E��@#������UH��H����H�����I��     L�H�}�H�}� t7H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@����H�E��P������UH��H��(��H�����I�)     L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H��(��H�����I��     L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H����H�����I�     L�H�}��E�_   �(�E�Hc�H�E�H�� < u�E�Hc�H�E�H��  �m��}� y����    ����UH��H����H�����I�     L�H�}�H�E�H�E�H�E�H�E��H�E�� </uH�E�H��H�E�H�E�H�E�� ��u�H�E�����UH��H��0  ��H�����I��     L�H������H������H������H�E�H������H�E�H������H�E��E�    �?H�E�� ��u�E�Hc�H�E�H��  �H�E�H�PH�U��U�Hc�H�U�H�� ��E��}�_~��E�    �-H�E�H�PH�U��H�E�H�PH�U�� 8�t�   ��E��}�_~͸    ����UH��SH�� ��H�����I��     L�H�}�H�u�H�E؋PH�E؋@ЉE�E�H�U����H�8      H�H�¾   H���������H��ЉE�}� t
�������   �E�    ��   �E�%�  ��H�8      ��H؋���uf�E�%�  ��H�8      ��H��������E�H�U����H�8      H�H�¾   H� �������H��ЉE�}� t������r�E��m�E�%�  =�  uE�E��E�H�U����H�8      H�H�¾   H���������H��ЉE�}� t�������E�H�E؋@$9E����������H�� []���UH��H����H�����I�>     L؉}��u�H�U�H�M�    ����UH��AWSH��0��H�����I�     Lۉ}�H�u�H�U�H�EȋPH�Eȋ@ЉE�H�Eȋ@ �E܉E�ЉE�   �    H�8      H�<I��H�hC������H����E�    �B�U�E�Љ�H�EЋ ��H�8      H��   H� �������H��ЉE��}� u�E�H�EȋP �E�9�w���H��0[A_]���UH��H����H�����I�     L�H�}�H�u�H�U��R��H�U����H�U�H��H��   I���������J� ������UH��AWSH��`��H�����I��     L�H�}�H�u�H�U�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H��������H���H�E�H�E�H�E�H�E�H��I��H�i$������H��ЉE�H�E��@,�E��9  H�E�H�E��H�E�� </uH�E��  H�E��H�E�H�E�� ��u׋U�H�E��@ H�M��	��H�M���H���������H��ЉE؃}� t#H�E�H��I��H���������H��и    ��   �E�    �f�E���Hc�H�E�H�H�E�H�E��@a��t5H�E��@b����@��t#H�E�H�U�H��H��H�E�������H��ЉE���E������}� t�E��}�?~����}� u+�}�?%H�EЋ@k�E�H�E��@ �E؉E�ЉE�m��	�E�    �
�}� �����H�E�H��I��H���������H��ЋE�H��`[A_]���UH��AWSH��P��H�����I��
     L�H�}�H�u�H�U��M�L�E�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H��������H���H�E�H�Eغ    �    H��I��H�hC������H��ЋU�H�E��@ H�M��	��H�M؉�H���������H��ЉE�}� t#H�E�H��I��H���������H��и������   �E�    �T�E���Hc�H�E�H�H�E�H�E��@a��t#H�E�H�U�H��H��H�E�������H��ЉE���E������}� t�E��}�?~����}� u:�}�?4�E���Hc�H�E�H�H�EȺ�   H��H��I��H��B������H�����E�����H�E�H��I��H���������H��ЋE�H��P[A_]���UH��AWSH��P��H�����I��     L�H�}�H�u�H�U�H�E���C  ��u
������	  H�E���C  ��@v/H��������H�<I�߸    H�2r������H��Ҹ������  H�E��PH�E��@ЉE�H�E���?  H�E��@ �ЋE�ЉE�    I��H��������H���H�E�H�Eغ    �    H��I��H�hC������H��ЋU�H�E��@ H�M��	��H�M؉�H���������H��ЉEԃ}� t!H�E�H��I��H���������H��ЋE��  H�E���C  ��H��H��H�E�H�H�E�H�EȺ`   �    H��I��H�hC������H���H�E�H��+H��H���������H���H��H�E�H��H��I��H��E������H����E�    �"H�UȋE�H����uH�UȋE�H�� �E��}�_~�H�E��@` H�E���+  H�EȉPo�U�H�E��@ H�M��	��H�M؉�H� �������H��ЉE�H�E�H��I��H���������H��ЋE�H��P[A_]���UH��AWSH��`��H�����I�     L�H�}�H�u�H�U��S  I��H��������H���H�E�H�EкS  �    H��I��H�hC������H���H�E��PH�E��@ ��H�EЉP�    I��H��������H���H�U�H�BH�E��PoH�EЉ�+  H�E��PH�EЉ�/  H�E��P H�EЉ�3  H�E��H�EЉ�G  �    I��H��������H���H�U�H��K  H�E�H��K  �    �    H��I��H�hC������H���H�E��@k�E�    I��H��������H���H�E��E������E�    �E�    ��  �   I��H��������H���H�U�H��K  �M�Hc�H��H�H�H�E�H��K  �U�Hc�H��H�H� H�E�H�E��   �    H��I��H�hC������H����E�    �<  H�E��@ �E��H�E��@�H�E��P�E�H�H�4�    H�E�H�ʉH�EЋ�;  �PH�EЉ�;  �E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E�;E�ts�E�H�U����H�U�H��H�¾   H���������H��ЉE��}� t:H�E�H��I��H���������H���H�E�H��H�o������H��и    �   �E��E�H�E��@�����E�    ��U�E�H��    H�E�HЋ �E�}��u	�E�������E��}��  ������}��t�E��}��  � �����H�E�H��I��H���������H���H�E�H��`[A_]���UH��AWSH��p  ��H�����I��     L�H������H�������   I��H��������H���H�E�H�E�H�E�H�E�H   H�E�H������H�E�H��H��I��H�&"������H���H�U�H�E�H��H��I��H��$������H��п�   I��H��������H���H�      H�H�      H���   �    H��I��H�hC������H��п   I��H��������H���H�E�H�EȺ   �    H��I��H�hC������H���H�E�H�E�H�E��   �    H��I��H�hC������H����E�    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ ���    Hǅ���    Hǅ���    Hǅ���    Hǅ ���    Hǅ(���    Hǅ0���    Hǅ8���    Hǅ@���    HǅH���    HǅP���    HǅX���    Hǅ`���    Hǅh���    Hǅp���    Hǅx���    H�E�    H�E�    H������H������H��H��I��H��E������H���������<wt������<au�E�   H�E��@   H�E��     H�U�H�E�H��H��H���������H��ЉE�}� t_H�      H�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��и    �  H�E�H�U�H�M�H�E�H��H��H�6�������H��ЉE��}� u_H�      H�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��и    �  H�EȋU��P,H�      H�H�M�H�U�H�u�I�ȹ    H��H�K�������H��ЉE�}����   �}� tqH�      H�H������H�U�H�u�A�    H��H�������H���H�      H�H������H�U�H�u�I�ȹ    H��H�K�������H��ЉE�}� ��   H�      H�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��и    ��  �}� t_H�E�H��I��H���������H���H�      H�H��I��H���������H���H�E�H��I��H���������H��и    �r  H�      H�H�U�H�M�H��H��H�r�������H���H�E�H�}� ��   H�      H�H��H�E�H��+�`   H��H��I��H��B������H���H�E�H��+H��H�u�������H���������<wt������<+t������<au
H�E��@"�H�E��@"H�E��@   H�EȋP,H�E���?  H�      H��PsH�E���C  ������<auH�      H��PoH�E��P#H�E�H��I��H���������H���H�      H�H��I��H���������H���H�E�H��I��H���������H���H�E�H��p  [A_]���UH��AWSH��@��H�����I���      L�H�}��   I��H��������H���H�E�H�E�   �    H��I��H�hC������H���H�E�H�E�H�E�   �    H��I��H�hC������H���H�E��@   H�E��     H�U�H�E�H��H��H���������H��ЉE܃}� t H�E�H��I��H���������H��и�����AH�U�H�M�H�E�H��H��H��������H��ЉE�H�E�H��I��H���������H��ЋE�H��@[A_]���UH��AWSH�� ��H�����I���      L�H�}�H�E�H�@H��I��H���������H����E�    �TH�E�H��K  �U�Hc�H��H�H� H��t?H�E�H��K  �U�Hc�H��H�H� H��I��H���������H��ЃE��}��  ~���H�E�H��K  H��I��H���������H���H�E�H��I��H���������H���H�E�    �    H�� [A_]���UH��H�� ��L�����I���      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H���������I� ������UH��H�� ��L�����I���      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H� �������I� ������UH��AWSH��   ��H�����I���      L�H��x���H��p�����l����   I��H��������H���H�E�H�E�H�E�H�E�H   H�E�H��x���H�E�H��H��I��H�&"������H���H�U�H�E�H��H��I��H��$������H��п   I��H��������H���H�E�H�EȺ   �    H��I��H�hC������H���H�E�H�E�H�E��   �    H��I��H�hC������H���H�E��@   H�E��     H�U�H�E�H��H��H���������H��ЉE��}� t_H�      H�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��и�����-  H�E�H�U�H�M�H�E�H��H��H�6�������H��ЉE��}� u_H�      H�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��и�����  H�EȋU��P,H�EȋPH�Eȋ@ЉE�H�EȋP,H�Eȋ@ �ЋE�ЉE��    I��H��������H���H�E�H�E��    �    H��I��H�hC������H��ЋU�H�Eȋ@ H�M��	��H�M���H���������H��ЉE��E�    �E�    �   �E���Hc�H�E�H�H�E��E�;�l���}~H�E��@a��ta�E���Hc�H��p���H�H�E���   H��H��I��H��B������H��ЋE���Hc�H��p���H�H��H�u�������H��ЃE����E��}�?�e�����H�E�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��ЋE�H�Đ   [A_]���UH��AWSH��`��H�����I���      L�H�}�H�u�H�U�H�M�D�E�H�E�H�E�H�Eغ�   �    H��I��H�hC������H���H�E�H��H���������H���H��H�E�H��H��I��H��E������H����E�    �"H�U؋E�H����uH�U؋E�H�� �E��}�_~�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉEп    I��H��������H���H�E�H�EȺ    �    H��I��H�hC������H��ЋU�H�E��@ H�M��	��H�Mȉ�H���������H��ЉEă}� t!H�E�H��I��H���������H��ЋE���  �E�    �$�E���Hc�H�E�H�H�E�H�E��@a��t�E��}�?~���H�E��@a���G  �}�?�=  �U�H�E؉PsH�E��@a��E���H�E؈PbH�U�H�E�H��H��H�,�������H���H�U؉BkH�E؋@k���uOH�E�H��H�,�������H�<I�߸    H�2r������H���H�E�H��I��H���������H��и   ��   �E���@��t$H�E؋@kH�U�H�M�H�Ή�H���������H���H�M�H�E຀   H��H��I��H��B������H��ЋU�H�E��@ H�M��	��H�Mȉ�H� �������H��ЉEĐH�E�H��I��H���������H��и    �JH�E�H��I��H���������H���H�E�H��H�P�������H�<I�߸    H�2r������H��Ҹ����H��`[A_]���UH��AWSH��P��H�����I���      Lۉ}�H�u�H�U��    I��H��������H���H�E��E�    �E��E��E������E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E��E܋E�;E���   �}� tV�E�H�U����H�U�H��H�¾   H� �������H��ЉẼ}� t#H�E�H��I��H���������H��и�����?  �E�H�U����H�U�H��H�¾   H���������H��ЉẼ}� t#H�E�H��I��H���������H��и������   �E��E�E��E��E�   H�E��@�����E�    ��U�E�EȋE�H��    H�E�HЋ �E�E�H��    H�E�H��     �}��uL�E�H�U����H�U�H��H�¾   H� �������H��ЉE̐H�E�H��I��H���������H��ЋE��6�E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��Y���H��P[A_]���UH��AWSH��   ��H�����I�7�      L�H��h����   I��H��������H���H�E�H�E�H�E�H�E�H   H�E�H��h���H�E�H��H��I��H�&"������H���H�U�H�E�H��H��I��H��$������H��п   I��H��������H���H�E�H�E��   �    H��I��H�hC������H���H��p���H�E�H�E��   �    H��I��H�hC������H���H�E��@   H�E��     H�U�H�E�H��H��H���������H��ЉE�}� t<H�E�H��I��H���������H���H�E�H��I��H���������H��и    ��  H�E�H�U�H�M�H�E�H��H��H�6�������H��ЉE��}� u<H�E�H��I��H���������H���H�E�H��I��H���������H��и�����d  H�E��U��P,H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE��    I��H��������H���H�E�H�E��    �    H��I��H�hC������H��ЋU�H�E��@ H�M��	��H�M���H���������H��ЉE�}� tSH�E�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��ЋE��l  �E�    �   �E������E���Hc�H�E�H�H�E�H�E��@a��t!H�E�H�U�H��H��H�E�������H��ЉE�}� u9H�E��@a �U�H�E��@ H�M��	��H�M���H� �������H��ЉE�}� ��E��}�?�k����}� tPH�E�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��ЋE��uH�E��@kH�U�H�M�H�Ή�H�o������H��ЉE�H�E�H��I��H���������H���H�E�H��I��H���������H���H�E�H��I��H���������H��ЋE�H�Đ   [A_]���UH��H����H�5����I���      Lމ}�E�E��}� u�E��   �E����rH�H     H�H�H     H�����UH��H����H�����I�w�      L�H�}��   H�E�H���r�����UH��AWH����H�����I�<�      L�H�8     H�H�U�H�@     H�    H���      �    H�M�   �    H��I��H�hC������H��ѐH��A_]���UH��AWSH��P��H�����I���      Lۉ}��u��}� u
�    ��  H�@     H�H=�   v%H���������H�<I�߸    H�2r������H��ҐH���      ���u�H���      ��PH���      ��E����E�E�%�  ��t�E��E�    �E�    �E�    �}� t�E��   �E�   �K  �}��  �=  H�8     H�H�E�H�E�    �E�    �  H�E؋@����   H�E؋@9E���   H�E�H�H�E؋@��H�H�E�H�E؋@+E���H�E؉PH�E؋P�E��H�E؉PH�E�H�E�H�8     H�H�E��E�    �mH�E؋@��tH�E��E��WH�E�H�E�H�E�H�E�H�E�H�@H�PH�E�H�PH�E��@   H�E�H�U�H�H�E��U��PH�E�H�U�H�P�E���!�}��   ~��H�E��E��}��   ������E�   ���}� ��   H�8     H�H�E��E�    �~H�E؋@��tH�E��E��hH�E�H�E��E��H�������H���H�E�H�E�H�U�H��E��E���H�E��PH�E��U��P�E���+E���H�E��PH�E�H�@   ��}��   �u���H���      �    H�@     H�H�PH�@     H�H�E�H��P[A_]���UH��SH��(��H�����I���      L�H�}�H�}� ��  �H���      ���u�H���      ��PH���      �H�E�H�E�H�8     H�H�E��E�    �M  H�E�H� H9E�tH�E��E��2  H�E�H�E�H�@     H�H�P�H�@     H�H�E؋@��uH�E�H��H�}������H����   H�E؋@��uH�E�H�@H�E�H�E�H�@H�P�H�E�H�PH�E�H�@H��tH�E؋@����   H�E�H�@H��uRH�E�H� H��H�}������H���H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    ��}��   �������H���      �    ��H��([]���UH��AWH��H��L�����I���      M�H�}��u�H�E�    �E�    H�}� u�E��   ��H�=������I� ���8  �H���      A� ��u�H���      A� �PH���      A� H�8     I� H�E�H�E�H�E��E�    �   H�E�H� H9E�t
H�E��   H�E�H�E��E�   H�E��P�E��=   v@H�@     I� �U�H�E�H��H���������I�< M�Ǹ    I�2r������M�A����H�E�H� H�E�H�E��P�E��H�E��P�E��}��   �X���H���      A�     �}� u�E��   ��H�=������I� ���H�E�H��HA_]���UH��H�� ��H�����I���      L�H�}�H�u��E�    H�E�H�E��   H�E�� ��H�E��@9�sH�E��P#H�E��@9�rH�E��@#    H�E�f�   H�E�H�PH�E��@#��H�H�E�H�PH�E�H�PH�U�H�U�H�R� �H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  �E��}��E����E�����UH��H�� ��H�����I���      L�H�}�H�u��E�    H�E�H�E�H�E��@'�PH�E��P'H�E��P'H�E��@9�rH�E��@'   �H�E��P#H�E��@'9�r�H�E��@'�P�H�E��P'�JH�E�H�PH�E��@'��H�H�E�H�PH�E�H�PH�E�H�HH�M���H�E��@'�PH�E��P'�E��}�~��E�����UH��AWSH��0��H�����I��      L�H�}�H���������H�H� H�E�H�E�H�E�H�E�H��I��H��H������H��ЉE�H�E�H��I��H��H������H��ЉE؋U܋E��=   ~
������   H�E�� </uH�E��E�H�HE�H�m�H�E�� </tH�E�H�E�H�PH�U�� /�H�E�H�U�H�E�H��H��I��H��E������H���H�E�H��I��H��H������H��Љ�HE�H�m�H�E�� </u	H�E��  �H�E�H�E��  �    H��0[A_]���UH��AWSH����H�����I���      L�H���������H�H� H��I��H��H������H��Ѓ�w
�    �   H���������H�H� H�E�H�E�H��I��H��H������H��Љ�HE��H�E�H�P�H�U��  H�E�� </u�H���������H�H� H��I��H��H������H��Ѓ�vH�E��  �    H��[A_]���UH��AWSH��0��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
�    ��  H�E�H��I��H��H������H��ЉE�E�H�H�P�H�E�H�� </u�E�H�H�P�H�E�H��  �}� 
�    �  �}���   H�E�H��� <:u%H�U�H�E�H��H��I��H��E������H����K  H��������H�<I��H�]�������H���H��H�E�H��H��I��H��E������H���H�E�H��I��H��H������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H��E������H����   H��������H�<I��H�]�������H���H��H�E�H��H��I��H��E������H���H�E�H��I��H��H������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H��E������H���H�E�H��0[A_]���UH��H����H�����I���      L�H�}�H�E�H�E�H�}� u�    �+�E�    �H�E�� </u�E�H�E�H�E�� ��u�E�����UH��AWSH��0��H�����I��      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
������   H�E�H��I��H��H������H��ЉE�E�H�HE�H�m��H�E�� </tH�m�H�E�� ��t�E�P��U�����H�E�H�U�H�E�H��H��I��H��E������H���H�E��  �    H��0[A_]���UH��H��0��H�����I�8�      L�H�}�H�u��U܉M�L�E�H���������H�H� H�E��E�H9E�}?H�E��@��H9E�}0H�E�H�E��E�H�E�H��H�E�H�H��    H�E�HE؉������UH��SH��@��H�����I���      Lۉ}ԉuЉỦM�L�E�L�M�f�E�  H�E�H�@H�E�H�E��@�E�}�u�E�    �E�    �   f�E� H�E��@�EȉE��H�H� H�E�H�� f�E�H�E�� ���E��J�E�f#E�f��t5�UЋE��Hc��UԋE��H�H�}��M�U�I��H��H��%������H���f�e�m��}� y��E�H�E��@9E��b�����H��@[]���UH��AWSH��0��H�����I���      Lۉ}܉u؉UԉM�D�E�L�M��E�    �X�E�    �CH�E�L��   �M�H�E��P�u؋E��Hc��}܋E��H�H��I��H��%������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I���      Lۉ}܉u؉UԉM�D�E�L�M��E�    �p�E�    �[H�E�H��   �E��E�i��E��A��H�E��P�M؋E��Hc��M܋E��H�I��D��H��I��H��%������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I��      Lۉ}܉u؉UԉM�D�E�L�M��}� �[  �}� �Q  �E�    �>H�E�L��   �M�H�E��P�E�Hc��}܋E��H�H��I��H��%������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E����Hc��}܋E��H�H��I��H��%������H��ЃE��E�;E�|��E�    �AH�E�H��   �M�H�E��P�u؋E��Hc��E�H�I��H��I��H��%������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E��Hc��}܋E����H�H��I��H��%������H��ЃE��E�;E�|���H��0[A_]���UH��AWSH��@��H�����I�j�      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}��  �E�    ��   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��   �E�f#E�f��tDH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H��%������H����BH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H��%������H���f�e�m��}� �[����E�H�E��@9E��	�����H��@[A_]���UH��SH��8��H�����I��      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H��*������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I�D�      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}���   �E�    �   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��W�E�f#E�f��tBH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H��%������H���f�e�m��}� y��E�H�E��@9E��T�����H��@[A_]���UH��SH��8��H�����I�'�      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H��,������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I�i�      L�H�}ȉuĉU��M�D�E�D�M�H���������H�H� H�E�H�E�H   � �? �    H��I��H�hC������H����E�    �U�H�E��P4�UH�E��P8�UH�E��P<H�E��@H   H�E��@L   H�E��P<H�E��PP�UH�E��PTH���������H�H��H�E�H�PXH�E��@D    H�E��PDH�E��P@�U�H�E��P�U�H�E��P�U�H�E��P �U�H�E��P�U H�E��P`�} u�E�   H�E��@�P�H�E��P(H�E��P�E�)ЍP�H�E��P$H�E��@0   �E����H�E��P,H�E��@��H�E��@��H�E�I���Ѻ    �    I��H�)?������H���H�E��@4��H�E��@����H�E�I��A�ȹ   �   �   H�g'������H��Ѓ}� u:H�E��@����H�E�I��A���� �   �   �   H�g'������H����8H�E��@����H�E�I��A���� �   �   �   H�g'������H��Ѓ}� t}H�E��@����H�U��E�I��A���� ����   �   H�g'������H���H�E��@4��H�E��@���ƋE��H�U�I��A�ȹ   ��ƿ   H�g'������H���H�E��@8A��H�E��@$��H�E��@(��H�E��@,��H�E��@0��H�E�I��H�g'������H���H�E�H��I��H��H������H������E�H�E�H�pHH�E��@��E܉������)Љ�H�E�H���u�I��A���� ������   ��H��H��-������H���H��H�E��@����H�E�I��A�    �   �   �   H��(������H���H�E�H�PHH�E��@��H���u�I��A���� ������   �ƿX   H��,������H���H��H�E�H�PHH�E��@��(H���u�I��A���� ������   �ƿ-   H��,������H���H��H�E�H�e�[A_]���UH��AWSH��0��H�����I���      L�H�}�H�u�H�E��P0H�E��@Ѓ�P�E�H�E��P,H�E��@Ѓ��E��E�P   �E�   �E�    �E���� H�E�H��I��H��H������H��ЉE�H�E�L�@H�M؋U܋E���������p��E�<�E��������ƋE���)ƋE��H�E�H���u�M��A�ȉщ�H��H��+������H���H���H�e�[A_]���UH��H����H�����I���      L�H�}��   H�E�H���r�����UH��H����H�����I���      L�H�}������UH��H����H�����I�}�      L�H�}�H�U��BD    H�U��JDH�U��J@H�U��R8A��H�U��R$��H�U��R(A��H�U��R,��H�U��R0��H�U�I��D��I�g'������J��А����UH��SH��(��L�����I���      Mډ�f�E�H���������I�H� H�E�H���������I�H��H�E�H�PXH�E�@(�P�H�E�@H���к    ��E�H�E�@$�P�H�E�@L���к    ��E�H�E�P<H�E�PPH�E�PD�E�9�rH�E��@D    H�E�@@�PH�E�P@H�E�P@�E�9�r9H�E��@D    H�E�PDH�E�P@H�E�H��H�w4������I����E��  f�}���   H�E�@D����   H�E�@D�P�H�E�PDH�E�H�xHH�E�pTH�E�@PH�U�J,H�U�RLA��H�U�R@A��ʃ���H�U�J0H�U�RHA��H�U�RDA��ʃ�A��H���u�I��A������D�޿    H��*������I���H����   f�}�	uH�E�@D�PH�E�PD��   f�}�
u!H�E��@D    H�E�@@�PH�E�P@�   f�}���   H�E�H�xHH�E�pTH�E�PPH�E�H,H�E�@LA��H�E�@@A��ȃ���H�E�H0H�E�@HA��H�E�@DA��ȃ�A���E�H���u�I��A���щ�D�މ�H��*������I���H��H�E�@D�PH�E�PD�E�H�]�����UH��H����H�����I�*�      L؉}�H���������H�H� H�E��U�H�E��P<�����UH��SH��(��H�����I���      L�H�}�H�}� t=H�E�H�E��&H�E�H�PH�U�� f�����H�5������H���H�E�� ��u���H��([]���UH��AWSH��P��H�����I�i�      L�H�}��u��U��M�L�E�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H��������H�<I�߸    H�2r������H��Ҹ�����6  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H��������H�<I�߸    H�2r������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�6�������H�<I�߸    H�2r������H��Ҹ   ��   �E�    �   �E�    �   �}� tNH�E�H��   H�E��P�M��E���E��Hc��M��E���E��H��M�I��H��I��H��%������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H��%������H��ЃE��}� �U����E��}� �;����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��P��H�����I���      L�H�}��u��U��M�D�E�L�M�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H��������H�<I�߸    H�2r������H��Ҹ�����3  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H��������H�<I�߸    H�2r������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�6�������H�<I�߸    H�2r������H��Ҹ   ��   �E�    �   �E�    �   �}� tKH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H��%������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H��%������H��ЃE��}� �X����E��}� �>����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��0��H�����I���      Lۉ}܉u؉U�H�M��E�    �   �E�    �t�U�������E��H�x�������H�Hڋ��E�}� tBH�E�H��   H�EȋP�MԋE��Hc��M؋E��H��M�I��H��I��H��%������H��ЃE��}�~��E��}��o�����H��0[A_]���UH��AWSH��@��H�����I���      Lۉ}̉uȉUĉM�L�E��E���� �E�``` �E���� �EĉE��ẺE܋E��E؋EȉEԋE؍P��E��xH�M��E�I��A�    �   ��I��H��(������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H��(������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H��(������H��ЋEԍP��E܍pH�M��E�I��A�    �Ѻ   ��I��H��(������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H��(������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H��(������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H��(������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H��(������H��ЋEԍP��E܍p�M��E�ȃ�H�M�I��A�    �Ѻ   ��I��H��(������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H��(������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H��(������H��ЋE؍P��M܋E�ȍp��E���H�M�I��A�    �   ��I��H��(������H��АH��@[A_]���UH��H��8��H�����I���      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �CH�E�H�PH�U�� ���E�H�E�H�PH�U�� ���E�E�+E�E�}� u�}� t
�m��}� u��E�����UH��H��8��H�����I��      L�H�}�H�uЉŰẺE�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M����E��P��U���u�H�E�����UH��H�� ��H�����I���      L�H�}���U��E�E��E�H�E�H�E��H�E�H�PH�U��U��m��}� u�H�E�����UH��AWSH��0��H�����I�'�      L�H�}�H�u�H�E�H�E�H�E�H�E��E�    H�E�H�PH�U�� ����I��H�
R������H��ЉE�H�E�H�PH�U�� ����I��H�
R������H��ЉEԋE�+EԉE܃}� u�}� t뗋E�H��0[A_]���UH��AWSH����H�����I�l�      L�H�}�H�u�H�E�H��I��H��H������H��Љ�H�E�H�H�E�H��H��I��H��E������H���H�E�H��[A_]���UH��H�� ��H�����I���      L�H�}�u�H�E�H�E��H�E�� ��9E�uH�E��H�E�H�E�� ��u۸    ����UH��H�� ��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E��3H�E��H�E�� 8�u!H�E�� ��H�E�� ��Ѕ�u�    �'H�E�H�PH�U��H�E�H�PH�U�� 8�t����������UH��H��0��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E��  H�E�����UH��AWH��(��H�����I�}�      L�H�}؉uԋU��҉Uԃ}� uOH�U�H��I��H��H������H��҉�H�E�H���   H�E�� ��tH�E�� ��9E�u	H�E��   H�E�H�E؃�H��űE�i��E�H�E�H�E��H�E�H�E� ������H�E� ��!�%������u%H�E� 3E䍐����H�E� 3E���!�%������t�H�E�H�E��H�E�H�E�� ��tH�E�� ��9E�u�H�E�H��(A_]���UH��H��@��H�����I�T�      L�H�}�H�u�H�U�H�U�H�U������   H�U�H�������   H�E�    H�E�    H�E�    H�E�    �H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�t�H�E�H+E��'H�U����H�Uȉ�H��H�uF������H���H+E�����UH��H����H�����I��      L�H�}�H�E�H�E��H�E�H�E�� ��u�H�E�H+E�����UH��AWSH��@��H�����I�϶      L�H�}�H�u��U�H�E�H�E�H�E�H�E��E�    �kH�E�H�PH�U�� ����I��H�
R������H��ЉE�H�E�H�PH�U�� ����I��H�
R������H��ЉEԋE�+EԉE܃}� u�}� t
�m��}� u��E�H��@[A_]���UH��H��(��H�����I�
�      L�H�}�H�u��U�H�E�H�E�H�E�H�E��}� u)������2H�E�H�PH�U��H�E�H�PH�U�� 8�u�m��}� u����E�����UH��H��8��H�����I���      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �!H�U�H�BH�E�H�E�H�HH�M����E��E�9E�w�H�E��  �E�����UH��AWH����H�����I��      L�H�}�H�u�H�M�H�U�H��H��I��H��G������H��҉�HE�H�E�� ��tH�E���    H��A_]���UH��AWH��(��H�����I���      L�H�}؉u�H�U�H��I��H��H������H��҉E��U�H�E�H�H�E��E�    �H�E�� ��9E�uH�E��H�m��E��E�9E�wڸ    H��(A_]���UH��H��0��H�����I��      L�H�}�H�u�H�E�H� H�E�H�}� u�    �vH�E�H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u,�}� u
H�E�    �H�E�H���  H�E�H�U�H�H�E���}� u������UH��H��@��H�����I�K�      L�H�}�H�u�H�E�H�E�H�E�    H�E�    H�E�    H�E�    H�E�� ��u
�    ��   H�E�H��� ��u+�H�E�H�E��H�E�� 8�t�H�E�H+E��   H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�u�H�E�H+E�����UH��H��8��H�����I��      L�H�}�H�u�H�U�H�}� uH�E�H� H�E�H�}� u
�    ��   �H�E�H�PH�U�� ���E�H�E�H�E��
�E�;E�u��H�E�H�PH�U�� ���E��}� uۃ}� uH�E�H�     �    �   H�E�H��H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u4�}� u
H�E�    �H�E�H��H�E�H�E��  H�E�H�U�H�H�E���}� u������UH��H����H�����I��      L�H�}�H�u�H�u�H�M�H���      H�H��H��M������H�������UH��AWSH�� ��H�����I���      L�H�}�H�u�H�E�H��I��H��H������H��ЉE��2�U�H�M�H�E�H��H��I��H�[B������H��Ѕ�uH�E��H�E�H�E�� ��uø    H�� [A_]���UH��AWSH�� ��H�����I��      L�H�}�H�E�H��I��H��H������H��Ѓ��E�E��I��H��������H���H�E�H�}� u�    �$�U�H�M�H�E�H��H��I��H��B������H��АH�� [A_]���UH��H��8��H�����I�R�      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��U�H�E�H�H�E�H�E�H;E�v[H�E�H;E�sQH�E�H�E��E�HE��H�m�H�m�H�E��H�E��H�E�H;E�u��'H�U�H�BH�E�H�E�H�HH�M���H�E�H;E�u�H�E�����UH��AWH����H�����I���      L�H�}�H�u�H�M�H�U�H��H��I��H�`E������H���H��A_]���UH��AWH����H�����I�8�      Lډ}�H�P�������H�<I�׸    H�2r������H�������UH��H����H�����I��      L؉}��U���H���������H�Hc��������t�E� �E�����UH��H����H�����I���      L؉}��U���H���������H�Hc��������t�m� �E�����UH��AWSH��0��H�����I�=�      L�H�}ȉuĉU��M��U�H�E�H��H�x�������H�<I�߸    I�2r������I�A��H�E�H��I��H���������H���H�E�H�E� �E�H�E� 9E�u��H��0[A_]���UH��AWSH�� ��H�����I���      L�H�}�H�u�H�E�� ��u�    �LH�E�� <wuH�E�H��I��H��X������H���H�U�H�E�H��H��I��H��������H���H�E�H�E�H�� [A_]���UH��AWH����H�����I��      L�H�}�H�U�H��I��H�q�������H���H��A_]���UH��AWH����H�����I���      L�H�}�H�U�H��I��H���������H���H��A_]���UH��AWH����H�����I�p�      L؉}�H�u�H�M��U�H�Ή�I��H���������H���H��A_]���UH��AWSH�� ��H�����I��      L�H�}�H�}� u������VH�E�H��I��H���������H��ЉE�H�E؋@��u+H�8�������H�H��E�H�։�I��H���������H��ЋE�H�� [A_]���UH��AWH����H�����I���      L؉}�H�u�H�M��U�H�Ή�I��H��T������H���H��A_]���UH��AWH����H�����I�2�      L�H�}�H�U�H��I��H��T������H���H��A_]���UH��AWSH��@��H�����I��      L�H�}ȉu�H�U�H�}� u	H�E��  H�E�H�E�H�E�H�E��E�    H�E�H��I��H���������H��ЉEԃ}����   H�E��@��u7�}�u�}� ~+H�8�������H�H��E�H�։�I��H���������H��Ѓ}�
tk�E�;E�}E�}�u�}� ~H�E�H;E�vH�m��m��:�}��^���H�E�H�PH�U�UԈ�E��D����}�u�}� ~�m���E��)�������}�~	H�E��  ��Eԉ�H�E�H�E�H��@[A_]���UH��AWSH�� ��H�����I���      L�H�}�H�u�H�}� u�    �^�E�    �2�E�Hc�H�E�H�� ��H�U�H�։�I��H��T������H��ЃE�H�E�H��I��H��H������H��ЋU�9�w��E�H�� [A_]���UH��AWH��(��H�����I��      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I���������I�A��H��(A_]���UH��AWH��(��H�����I���      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I���������I�A��H��(A_]���UH��AWH����H�����I�.�      L�H�}�H�U�H��I��H��������H���H��A_]���UH��AWH����H�����I��      L�H�}�H�U�H��I��H�b�������H��ҐH��A_]���UH��AWH��(��H�����I���      L�H�}�H�u��U܋U�H�u�H�M�H��I��H�C�������H���H��(A_]���UH��H����H�����I�@�      L�H�}�H�}� u������!H�E��P#H�E���+  9�r�������    ����UH��AWH����H�����I��      L�H�}�H�U�H��I��H�!�������H���H��A_]���UH��AWSH��`  ��H�����I���      L�H������H������H�������E�    �E�    �  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H��b������H���	E�}���  �E�H��    H�Q�  H�H�F�  H�>��H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E��E�H������H�։�I��H�mU������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�}� t(H������H�E�H��H��I��H�fW������H����O  H������H��H���������H�<I��H�fW������H����   H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E�H�������E�H�։�I��H�+�������H���H������H������H��H��I��H�fW������H����w  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������
   H��H��I��H���������H���H������H������H��H��I��H�fW������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������   H��H��I��H�r�������H���H������H������H��H��I��H�fW������H����  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�EȾ   H��fHn�I��H�`�������H���H������H������H��H��I��H�fW������H����]  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eк
   H��H��I��H���������H���H������H������H��H��I��H�fW������H����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ
   H��H��I��H���������H���H������H������H��H��I��H�fW������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ   H��H��I��H���������H���H������H������H��H��I��H�fW������H����G  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�E�   H��fHn�I��H�`�������H���H������H������H��H��I��H�fW������H����   H������H�ƿ%   I��H�mU������H��ЋE�Hc�H������H�� ��H������H�։�I��H�mU������H����4�E�Hc�H������H�� ��H������H�։�I��H�mU������H��ЃE��E�Hc�H������H�� ��������    H��`  [A_]���UH��H����H�����I��      L؉��E��E�    �E��S��%wa��H��    H�"�  H�H��  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I�\�      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H�XZ������L��Љ�<�����<���H���   A_]���UH��H�� ��H�����I�v�      L�H�}�H�u�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E�����UH��AWSH��  ��H�����I��      L�H������H������H��x����E�    H������H�E�f�E�  �E� �E�    �/  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H��m������H���	E܃}���  �E�H��    H���  H�H���  H�>��H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E��E�H�U�H�E�H��H��H�~d������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H�}� t'H�U�H�E�H��H��H�~d������H���H�E��e  H�E�H���������H�4H��H�~d������H���H�E��7  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E�H�������E�H�։�I��H�+�������H���H������H�E�H��H��H�~d������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������
   H��H��I��H���������H���H������H�E�H��H��H�~d������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������   H��H��I��H�r�������H���H������H�E�H��H��H�~d������H���H�E��3  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�E��   H��fHn�I��H�`�������H���H������H�E�H��H��H�~d������H���H�E��x  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�E��
   H��H��I��H���������H���H������H�E�H��H��H�~d������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ
   H��H��I��H���������H���H������H�E�H��H��H�~d������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ   H��H��I��H���������H���H������H�E�H��H��H�~d������H���H�E��e  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�Eо   H��fHn�I��H�`�������H���H������H�E�H��H��H�~d������H���H�E��   H�E�H���������H�4H��H�~d������H���H�E�fǅ����  �E�Hc�H������H�� ������H������H�E�H��H��H�~d������H���H�E��8�E�Hc�H������H�� �E�H�U�H�E�H��H��H�~d������H���H�E��E��E�Hc�H������H�� �������H�E��  H�U�H������H)�H��H�Ā  [A_]���UH��H����H�����I�5�      L؉��E��E�    �E��S��%wa��H��    H�L�  H�H�A�  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I���      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H��d������L��Љ�<�����<���Hc�H�����H��  ��<���H���   A_]���UH��AWH���   ��L�����I���      M�H����������H�����H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H����������H�����H��M��H�Wp������L��Љ�<�����<���H���   A_]���UH��AWSH��0��H�����I���      L�H�}؉u�H�U�H�M��}�   v
�    �   H�U�H�E�H��H���      H�<I��H��d������H��ЉE�}���  ~�   �I�E�E�}� ~:�U�H�E�H���      H�4H��I��H��B������H��ЋE�Hc�H�E�H��  �E�H��0[A_]���UH��AWH����H�����I�      L؉}�H�8�������H�H�
�U�H�Ή�I��H��T������H���H��A_]���UH��AWSH�� ��H�����I�e�      L�H�}�H�}� tj�E�    �?H�8�������H�H��E�Hc�H�E�H�� ��H�։�I��H��T������H��ЃE�H�E�H��I��H��H������H��ЋU�9�w���H�� [A_]���UH��AWH���   ��L�����I���      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�8�������I�H� H�� ���H�����H��H��M��H�XZ������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I�Ȍ      M�H��8���H��0���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�H���������I�<M�׸    H�2r������L�������UH��AWH����H�����I�*�      L�H�}�H�U�H��I��H��q������H��ҐH��A_]���UH��AWH��(��H�����I�ދ      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H�V������H��Ѹ    H��(A_]���UH��AWH��(��H�����I�y�      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H�V������H����H�E�H�E�� < tH�E�H   H9E�sH�E�� <
u�H�E��  H�E�H;E�����H��(A_]���UH��AWSH��0��H�����I�֊      L�H�}�H�uЉỦM�H���     H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H�V������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H���     H�H�E�H���     �0H���     �D �}�u-�U�H�E�    H��I��H�ڋ������H���H�U�H��   �}�u+�U�H�E�    H��I��H���������H��Љ�H�EЉ�[�}�u,�U�H�E�    H��I��H���������H��Љ�H�E�f��)�U�H�E�    H��I��H���������H��Љ�H�EЈ�    H��0[A_]���UH��AWSH��0��H�����I�2�      L�H�}�H�uЉỦM�H���     H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H�V������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H���     H�H�E�H���     �0H���     �D �}�u'H�E�H��I��H�K�������H����Z�H�E�� �+�}�u%H�E�H��I��H�K�������H���fH~�H�U�H��    H��0[A_]���UH��SH��8��H�����I���      L�H�}�H�u�H�U��E�    �E�    ��  �E�    �E�Hc�H�E�H�� ������%��  �E��E�Hc�H�E�H�� ������lu�E��E�   �E�Hc�H�E�H�� ����H�X|������H���	E�}��o  �E�H��    H��}  H�H��}  H�>��H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H�t������H�����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H�yt������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�u������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�u������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��v������H����?  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�u������H�����   H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�u������H����jH�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��v������H������E��E�Hc�H�E�H�� ��������E�H��8[]���UH��H����H�����I���      L؉��E��E�    �E��S��%wa��H��    H��z  H�H��z  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H��w������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I��      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H��w������L��Љ�<�����<���H���   A_]���UH��H����H�����I��      L؉}�H�u�H�}� u������w�}��u������jH�E��@#��tH�E��@#�P�H�E��P#H�E��@#H�U��J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U���E�����UH��AWSH����H�����I�]�      L�H���������H�H� H��I��H���������H��ЉE�}��t+H�8�������H�H��E�H�։�I��H���������H��ЋE�H��[A_]���UH��AWH��(��H�����I��      L�H�}�H�u�H�U�H���������H�<I�ϸ    H�2r������H�������UH��H����H�����I�z      L�H�}��	   H�E�H���r�����UH��SH����H�����I�@      L�H�}�H�}� u.H���     H�<H�z�������H���H���     H��H�E�H��H�z�������H���H�E�H��[]���UH��AWSH��0��H�����I��~      L�H�}�H�u�H�E�H���������H�4H��I��H�VS������H���H�E�H�}� u
������   �E�    H�E�H��I��H��H������H��ЉE܃}�`~	�E�   �$H�E�H�P+H�E�H��H��I��H��E������H���H�E��@���H�E��PH�E�H��I��H��S������H��ЋE�H��0[A_]���UH��H��0��H�����I��}      L؉}�H�u�H�E�H�E��E܉E��E�    �}� y,H�E�H�PH�U�� -�}�   �u�E�����E���E��؉E�H�E�H�E�M�Hc�Hi�gfffH�� ��������)�����)��ʉЍH0H�E�H�PH�U�ʈ�E�Hc�Hi�gfffH�� ����)ЉE�}� u��}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWSH��@��H�����I�|      L�H�}�H�u��U�H�}� u#H�E�H�E�H�E�H�PH�U�� 0H�E��  �  H�E�H�E؋E�Hc�H�E�H�H�E��3H�E؃��E�H�m��}�	~�7   ��0   �U��H�m���H�E�H�E�H;E�wËE�Hc�H�E�H��  H�E�H�E��E�    �8H�E�� <0uH�E��"H�U�H�E�H��H��I��H��E������H�����E��E�;E�|�H�E�H�E�H�E�H��I��H��H������H��Љ�H�E؋E�H�U�)Љ�H�M�H�E�HȾ    H��I��H�hC������H���H��@[A_]���UH��AWH����H�����I�{      L؉}�U�    ��I��H�=������H���H��A_]���UH��AWH����H�����I��z      L؉}�u�U��U��I��H��������H���H��A_]���UH��AWH����H�����I�oz      L�H�}�H�U�H��I��H�d������H��ҐH��A_]���UH��AWH����H�����I�#z      L�H�}�u�M�H�U��H��I��H�e������H���H��A_]���UH��H����H�����I��y      L؉}�u�E��}�E��E��}�ЉE��}� x�E���y�E����E��E�+E�E��!�}� y�E���~�E����E��U��E�ЉE�H�E�����UH��H�� ��H�����I�Jy      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H�� ��H�����I��x      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H��H��H�����I��w      L�H�}�H�u��U�H�E�H�E�H�E�H�PH�U�� ���E�E���H���������H�H������ ��uǃ}�-u�E�   H�E�H�PH�U�� ���E��"�E�    �}�+uH�E�H�PH�U�� ���E�}� t�}�u9�}�0u3H�E�� <xtH�E�� <XuH�E�H��� ���E�H�E��E�   �}� u�}�0u�   ��
   �E��}� t	H��   ������H�E�E�Hc�H�E�H�H��H�ЉE؋E�Hc�H�E�H�H��H�E�}� t�}� ~�E�)E�H�E��]�H�E�    �E�    �E���H���������H�H��������t�m�0�[�E���H���������H�H���������5  �E���H���������H�H��������t�7   ��W   )E�E�;E���   �}� ��   �}� tgH�E�H;E�|H�E�H;E�u0�E�;E�~(�E�����H�E�   �H�h�������H�� �����   �E�   �E�H�H�U�H��H�E��E�H�H)E��eH�E�H;E�H�E�H;E�u-�E�;E�~%�E�����H�E����H�h�������H�� �����$�E�   �E�H�H�U�H��H�E��E�H�HE���H�E�H�PH�U�� ���E��y������H�}� t�}� t
H�E�H���H�E�H�U�H�H�E�����UH��AWH����H�����I��t      L�H�}�H�M�
   �    H��I��H���������H���H��A_]���UH��AWH����H�����I�mt      L�H�}�H�M�
   �    H��I��H���������H���H��A_]���UH��AWAVAUATSH����H�����I�t      L�H�}�H�uȉU�L�eп    L��L�`� �؉���H���������H�H������ ��uЃ�-u�   L��L�`� �����+uL��L�`� �؃}� t�}�u-��0u(A�$<xt	A�$<XuI�D$� ��I���E�   �}� u��0u�   ��
   �EċE�Hc������    H��I�ǋE�Hc������    H��H�Љ�A�    A�    ����H���������H�H��������t��0�T����H���������H�H��������tz����H���������H�H��������t�7   ��W   )�;]�}GE��x
M9�wM9�u��9�~A������A�   �E�H�L��Hc�I�L��L�`� ���;������E��yA�����H�h�������H�� "   �	����tI��H�}� tE��tI�D$��H�E�H�U�H�L��H��[A\A]A^A_]���UH��H����H�����I��q      L؉}��   �   ���r����UH��AWSH����H�����I��q      L�H�}�H�E�H���������H�4H��I��H�`E������H��Ѕ�uH���������H�H� ��    H��[A_]���UH��AUATSH�� ��H�����I�q      L�H�}�H�u�H� �     ��E�L�e�H�]�E�,$L��L�`��H��H�XD�(�m��}� uې�H�� [A\A]]���UH��H��8��H�����I��p      L�H�}�H�u�H�U�H� �     ��E�H�E�H�E�H�E�H�E�H�E�H�E�H�E�� ���E�H�E�H�PH�U�H�U���H�E�H�PH�U�H�U���H�E�H�PH�U��U���m��}� u�������UH��SH��H��H�����I��o      L�H�}�H�u�H� �     ��E�H�E�H+E��EȋE�9E���  �E�����EȺ    ��E��EȋU�H�E�H�H�E�H�E�H�E�H�E�H�E�E�H�H��H��H�E�H�H�E�H�E�H;E�sjH��     H�H�U�H�E�H��H���щEă}� u/�E�H�H��HE�H�U�H�E�H��H��H�Ԏ������H�����  �}� y�E�H�HE���  �H�E�H;E���   H��     H�H�U�H�E�H��H���щEă}� u)�E�H�HE�H�U�H�E�H��H��H�Ԏ������H���뢃}� ��   H�E�H;E�uA�E�H�HE�H�U�H�M�H�E�H��H��H�O�������H��ЋE�H�HE�H�E�H�E��M���H�U�H�E�H��H��H�Ԏ������H��ЋE�H�H��HE��E�H�HE���   �E�H�H��HE�����H�E�H;E���   H�E�H+E�H��H�E�H+E�H9�|4�E�Hc�H�E�H�H�E�H��H��H���������H���H�E�H�E������H�U�H�E�H��H��H���������H��ЋE�Hc�H�E�H�H�E������E�H�H��HE�H�U�H�M�H�E�H��H��H�O�������H��ЋE�H�H��HE�H�E�H�E������H��H[]���UH��H�� ��H�����I�m      L�H�}��u�U�H�M�H��     H�U�H��U�H� �     ��U��U���H�U�H�H�U�H��H��H���������H��А����UH��AWH����H�����I��l      L�H�}�H���������H�<I�׸    H�2r������H��Ѹ����H��A_]���UH��H��@��H�����I�(l      L�H�}�H�u�H�U�H�U��H�E�H�U����H���������H�Hc���҃� ��u��E�    H�U���҃�+t��-u�E�   H�E�H�����������E��E�    �E�    �E�    �;�M�H�����������Y�H�U���҃�0�*��X��E�H�E��E�H�U����H���������H�Hc���҃���u�H�U����.uuH�E��?�M�H�����������Y�H�U���҃�0�*��X��E�H�E��E��E�H�U����H���������H�Hc���҃���u��U�)U�}� uH���������f���  �}� t�E�H���������f(fW��E�H�U����etH�U����E��   �E�    H�E�H�U���҃�+t��-u�E�   H�E��E�    �%�M܉����҉�H�U���҃�0ʉU�H�E�H�U����H���������H�Hc���҃���u��}� t�U�)U���U�U�}����|	�}�   ~H�����������   H�����������E��E�E܃}� yF�]��A�E܃���t&�}� y�E��^E��E���E��YE��E��}��E��Y��E��}� u�H�}� tH�E�H�U�H��E�����UH��H����H�����I��h      L؉}�H�E�   �E�    �H�U�H��H��H�H�H�E��E��E�;E�|�H�E�����UH��AWSH��@��H�����I��h      L��E�H�}��u�H�}� u	H�E��  H�E�H�E�H���������f��f/E�v,H�E�H�PH�U�� -�E�H���������f(fW��E��E�H��������f/s�E��H,�H�E��/�E�H����������\��H,�H�E�H�       �H1E�H�E�H�E�H�E�H��x�H*��H��H���H	��H*��X��M��\�f(��EȋE���H��������H���H��x�H*��H��H���H	��H*��X��YE�H��������f/s�H,�H�E��*H����������\��H,�H�E�H�       �H1E�H�E�H�E�H�M�H�U�H�E�H���������H�43H��I�߸    I�in������I�A��H�E�H��@[A_]���UH��AWH����H�����I��f      L�H�}�H�U�    H��I��H�̓������H���H��A_]���UH��AWH����H�����I�Wf      L�H�}�H�u�H�M�H�U�H��H��I��H�̓������H����Z�H��A_]���UH��AWH��(��H�����I��e      L�H�}�H�u�H�M�H�U�H��H��I��H�̓������H����E��E�H��(A_]���UH��H����H�����I��e      L؉}��E����3E�)�����UH��H��@��H�����I�me      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�    H�}� y>H�E�H�PH�U�� -H�       �H9E�uH��������H�E�H�E��H�E�H��H�E�H�E�H�E�H�M�H�gfffffffH��H��H��H��H��?H)�H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U��ʈH�M�H�gfffffffH��H��H��H��H��?H)�H��H�E�H�}� u�H�}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U߈H�E�H;E�w�H�E�����UH��AWH��8��H�����I��c      L�H�}�H�uЉU�H�U�H�U�H�}� yH�U�H�JH�M��-H�]�H�U�H�U��}�u$H�M�H�u�   H��I��H�r�������H����H�M�H�U�H��H��H���������H���H�E�H��8A_]���UH��H��0��H�����I�Hc      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E�H�M�H���������H��H��H��H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U�ʈH�E�H���������H��H��H��H�E�H�}� u�H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWH��8��H�����I�Mb      L�H�}�H�uЉU�H�U�H�U�H�U�H�U��}�u$H�u�H�M�   H��I��H�r�������H����H�M�H�U�H��H��H���������H���H�E�H��8A_]���UH��H����H�����I��a      L؉}������UH����H�����I��a      Lظ   ]���UH��H����H�����I�ia      L�H�}��    ����UH��H����H�����I�:a      L�H�}�H�`�������H�H� ����UH��H����H�����I��`      L�H�}�H�`�������H�H� ����UH��H�� ��H�����I��`      L�H�}��u�H�U�H�M�    ����UH����H�����I��`      Lظ    ]���UH��H����H�����I�c`      L��E�H��������f������UH��H����H�����I�*`      L��E�H��������f������UH��H����H�����I��_      L��E��}�H��������f������UH��H����H�����I��_      L��E�H�}�H��������f������UH��H����H�����I�x_      L��E��M�H��������f������UH��H��(��H�����I�:_      L��E��M��E��U��U��E��E��E������������������������������]��E�����UH��H����H�����I��^      L��E����E����]��E�����UH��H����H�����I��^      L��E�H��������f������UH��H����H�����I�X^      L��E�H� �������f������UH��H����H�����I�^      L��E�H�(�������f������UH��H����H�����I��]      L��E�H�0���������E��E�����UH��H����H�����I��]      L��E�H�8�������f������UH��H����H�����I�i]      L��E�H�@�������f������UH��H����H�����I�0]      L��E�H�H�������f������UH��H����H�����I��\      L��E�H�P�������f������UH��AWH����H�����I��\      L��E��E�H�X�������H�f(�fHn�I��H���������H���H��A_]���UH��H����H�����I�]\      L؉}�H�u�    ����UH��AWH����H�����I�)\      Lډ}�H�u�H�`�������H�<I�׸    H�2r������H�������UH��AWH��(��H�����I��[      Lى}�H�u�H�U�H�q�������H�<I�ϸ    H�2r������H�������UH��AWSH�� ��H�����I�|[      L�H�}�H���������H�<I�߸    H�2r������H����E�    �.�E�H�H��    H�E�HЋ ��I��H�0q������H��ЃE��}�?~̸����H�� [A_]���UH��AWH����H�����I��Z      L�H�}�u�H���������H�<I�׸    H�2r������H�����f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     fD                                                    "          "              "       "       "       "          "       "       "       !   "       !   "       !   "       !   "       !   "       !   "       !   "       !   "       !   "       !   "       !   "       !   "       !   "       "       "                                                                             !       !          !       !       !       !          !       !       !       !          !       !       !       !       !                                  !       !          !       !       !          !          !       !       !       !       !       !               	   !       !       !       !       !          !       !       !                  !       !             !       !       !          !          !       
   !       !          !          !              !          !                                                                                                	  
!           '(8    	                                        4/5*?7*+,-.03162,@-A.B90C1D2E4F5H:6I4G	"	#	#	#	#	#	#	#	#	#	#
$7J
%
%
%
%
%
%
%
%
%
%9K:L@PBQCRFSGTHUIVJW
&
&&=
&&=KXLY&>&>&>&>&>&>&>&>&>&>P\Q]))))))))))R^S_T`
&
&Va
&))))))))))))))))))))))))))WbXc<O<O)<O))))))))))))))))))))))))))!!Yd<O<O\e<O]f_g!!! `hcidjfkjlkm####################ln            !!    #;#;!!#;    !!        !!        $<$<$<$<$<$<$<$<$<$<    !!    !!#;#;  #;$&$&;M$&;M    ;N;N;N;N;N;N;N;N;N;N=>=>=>=>=>=>=>=>=>=>          $&$&  $&MNMNMNMNMNMNMNMNMNMNOZ  OZ    O[O[O[O[O[O[O[O[O[O[Z[Z[Z[Z[Z[Z[Z[Z[Z[Z[                 	
	"'++0000000000AAADDADAAAAAAAAAAAAAAAAAAAAAAADDADAAAAAAAAAAAAAAAAAAA                @(#)ncform 1.6 88/02/08 SMI    
   :<        ����       ��������   ����   (   A   [   _   .   a   ����\   ����   (   A   [   _   .   a   ����3   ����F     !     !   =   !     !   >   !   <   !     !     !     !   +   !   -   !   *   !   /   !   ����D   ����G   [   _   .   a   ����]   ����f             	     
          ����   ����u   ]   U   ����W   ����z        ����   �����     !     !   =   !     !   >   !   <   !     !     !     !   +   !   -   !   *   !   /   !   ����F   6   4   �   5      7   6   4      5      7      �         �      /   .   0   k   h   a   /   .   0   6   4   P   5      7   6   4   (   5   	   7   6   4   �   5   �   7   /   .   0   �   e   Q   /   .   0   
   6   4   ~   5   C   7   6   4   <   5   �   7   �   �   �   �   l   �   /   .   0   I      K   /   .   0         &   �      �      u   =   >   J      L   6         A   B   7   %   �   �   g   o   H      ]   ^   R   S   T   U   V   W   X   Y   Z   [   \   t   ;   M   6   4   v   5   c   7   n   _   @   ,   F   m      !   i   j   *   p   )   �   �         �   O   {   +   w      r   q   b   ?   �   �   z   D   '   $   �   #   x         f   }   �   �   N   E   F   G   �   �   �   �      |            y   `   �   �   �   �   �   �   s                                     �                   �                   �               �       �   �   �   �       �               �   �   �   �   �   9   :   1   2   3   8   9   :   1   2   3   8   �           d       -                   F                   9   :   1   2   3   8   9   :   1   2   3   8                       8                                           9   :   1   2   3   8           1   2   3   8                                                                    "           ����������������������"   ���������������+   ������(   ���������������]   �������+   +   +   \   ���������������+   +   ���+   ���>      ����0   S   ������+   +   +   +   +   +   +   +   +   +   +   ������Z      ���������+      ����(������<   ���������������+   ���+   Y   =   ������������������������������5   5   ������R   ����������������U      ���+   ������   +   �������8   <   ���������+   +   ����������������   "   ���+   ���   ������������?���      ����;   ����������:   +   ������������������&���!������+   �������   ���������   ���+   ����������������+   +   ���"   ���   ������������?������    �   2   `   G   �   �   �   �   �   �   �   �   �   �   R   6   �   �   �   �   �   ;   �   �   �   ?   F   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   E   �   �   A   �   �   �   L   �                                                                                                  !      "   #   "                                                   $                           &      '      %   %   )      (            *            +   +                     	   	   -   ,   
   
   .      0      /            1      2            3   4   3                                             	                                                                              	          	                                                      	   	                                                            	                                           	                  	                        	      	                                           �������������������    ��������  ����;   ����      ��������  ��������  ������������(   +   -   @   ����      ����  ��������=   ,   ����  ������������(     =   <   >         +   -   *   /         ��������������������(   ����������������������������,   ����=   [   .   (   ��������  ��������������������������������������������������������)   ����  ��������  	  ����,     ��������  ��������)   ,   ����������������{   [   )   ����������������������������]   )   ����  ������������������������  ��������������������������������������������    }   ,   ����]   ,   ������������  
  
  ������������=   ����
  ����  ����������������������������   ����             h                                           ����?   ^           !               0   ����4   5   6   7                         e               G                                                           !       .   /   K   =   8           	      ��������    c   f           B       H   I      #   $   %   &   '   (   )   *   +   ,   -   9   ;   "       L       >           ����E   e           b       C                      1   O   ����2             ����    d   g   `   @      J      :   <       P   Q   S       V              
          ����               M           N   Y   X   [       B                R                     T   Z                                                       ~ � � � � � � � � ~             ~ � � � � � � � � ~                 l � � � � | 8                   8 | � | 8                   < < � � �   <                < ~ � � ~   <                      < <              � � � � � � � � � � � � � � � �           < f B B f <           � � � � � � � � � � � � � � � �        2 x � � � � x             < f f f f <  ~               ? 3 ? 0 0 0 0 p � �              c  c c c c g � � �               � < � < �             � � � � � � � � � � �               > � >                  < ~    ~ <                f f f f f f f   f f              � � � {                | � ` 8 l � � l 8  � |                       � � � �              < ~    ~ <  ~              < ~                           ~ <                      �                         0 ` � ` 0                         � � � �                       ( l � l (                      8 8 | | � �                   � � | | 8 8                                                 < < <                  f f f $                             l l � l l l � l l           | � � � |   � � |               � �   0 ` � �             8 l l 8 v � � � � v           0 0 0 `                             0 0 0 0 0 0               0         0                   f < � < f                         ~                                    0                     �                                                           0 ` � �             8 l � � � � � � l 8              8 x       ~             | �    0 ` � � �             | �   <    � |               < l � �                 � � � � �    � |             8 ` � � � � � � � |             � �     0 0 0 0             | � � � | � � � � |             | � � � ~     x                                                       0                  0 ` 0                      ~     ~                     ` 0      0 `             | � �                       | � � � � � � � |              8 l � � � � � � �             � f f f | f f f f �             < f � � � � � � f <             � l f f f f f f l �             � f b h x h ` b f �             � f b h x h ` ` ` �             < f � � � � � � f :             � � � � � � � � � �             <         <                   � � � x             � f f l x x l f f �             � ` ` ` ` ` ` b f �             � � � � � � � � � �             � � � � � � � � � �             | � � � � � � � � |             � f f f | ` ` ` ` �             | � � � � � � � � |           � f f f | l f f f �             | � � ` 8   � � |             ~ ~ Z       <             � � � � � � � � � |             � � � � � � � l 8              � � � � � � � � � l             � � l | 8 8 | l � �             f f f f <     <             � � �   0 ` � � �             < 0 0 0 0 0 0 0 0 <               � � � p 8                 <         <          8 l �                                                   �       0                                     x  | � � � v             � ` ` x l f f f f |                   | � � � � � |                < l � � � � v                   | � � � � � |              6 2 0 x 0 0 0 0 x                   v � � � � � |  � x       � ` ` l v f f f f �                 8      <                        f f <       � ` ` f l x x l f �             8         <                   � � � � � � �                   � f f f f f f                   | � � � � � |                   � f f f f f | ` ` �             v � � � � � |                � v f ` ` ` �                   | � ` 8  � |              0 0 � 0 0 0 0 6                    � � � � � � v                   � � � � � l 8                   � � � � � � l                   � l 8 8 8 l �                   � � � � � � ~   �             � �  0 ` � �                 p                                        p         p                       v �                        8 l � � � �                               ��� ��� ~~~                                 uuu ��� ��� ���                                 ��� ��� ��� ��� ;;;                          ��� ��� ~~~ ��� ���                         ��� ��� ���     ��� ���                         ��� ���      ��� ��� ppp                 @@@ ��� ���         III ��� ���                 ��� ��� ��� ��� ��� ��� ��� ���                 ��� ���                 zzz ��� ���         ``` ��� ���                     ��� ���         ��� ��� MMM                     ��� ��� bbb     ��� ���                         ||| ��� ���      ��Cunexpected type to index table not enough memory        too few arguments to function `next'    too many arguments to function `next'   first argument of function `next' is not a table        error in function 'next': reference not found   r String: %10.10s... lua: %s
 function stack overflow   
	in statement begining at line %d in function "%s" of file "%s" 
	active stack
        	-> function "%s" of file "%s"
 
	in statement begining at line %d of file "%s" bad switch yylook %d    �I������VG�������I������G�������G�������G�������I�������G�������G�������G������H������H������H������H������)H������3H������=H������kH������uH������H�������H�������H�������H�������H�������H�������H�������H�������H�������H�������H������I������I������I������I������VI�������I������not enough memory       unexpected type at conversion to number string to number convertion failed      unexpected type at conversion to string %d %g   indexed expression not a table  internal error - table expected stack overflow  call expression not a function  internal error - opcode didn't match    "x�������U�������U������2V������V�������V������&W������}W�������W������KX�������X�������X������Y������RY�������Y�������Y������Z������ZZ�������Z�������Z������K[�������[�������\�������\������]������f]�������]������^������_^�������^������_������X_�������_������`������W`�������`������>a������%b������uc������?d�������d������ef������i�������j������&l������m�������m�������n�������o�������p������ q������^q�������q�������q������r������+r�������r�������r������s������v������Xw������bw�������w�������w�������f������e������;e������f�������e�������e������f������Bf������%g
 %s
 cfunction: %p
 userdata: %p
 table: %p
 nil
 invalid value to print
          �?   @  �B   �            type tonumber next nextvar print mark nil number string table function cfunction symbol table overflow not enough memory        lua: constant string table overflow string table overflow indexed table overflow too many files too few arguments to function `nextvar' too many arguments to function `nextvar'        incorrect argument to function `nextvar'        name not found in function `nextvar'    code buffer overflow stack overflow     too many local variables or expression too complicate variable buffer overflow  %s near "%s" at line %d in file "%s" out of memory yacc stack overflow syntax error     ¤������¤������3�������~�������¤������¤���������������������|�������¤������¤��������������¤������¤������¤������z�������6�������W�������Ʊ���������������������������¤������¤������¤�������������س���������������������¤������a�������ʹ������3���������������ֵ�������������7��������������ܶ������9���������������޷������&�������n�����������������������F�������\�����������������������@�������k���������������ƻ������0�������k���������������������J���������������ν�������������¤������E�����������������������־���������������������������^�������¤������¤������t�����������������������������"�������;�������T�������j�������������������������������G�������~����������������������������������������������#�������Z���������������%���������������������������������������x������������������������������¤������%�������  �?    c       usage: lua filename [functionnames] callfunc execstr test       incorrect argument to function 'readfrom` r     incorrect argument to function 'writeto` w %[^"]" %[^']' %s %%%ds %ld %f %% - %d .%d %c  
 %g   incorrect format to function `write'    incorrect argument to function 'execute` readfrom writeto read write execute remove   �?        too few arguments to function `abs'     incorrect arguments to function `abs'   too few arguments to function `sin'     incorrect arguments to function `sin'   too few arguments to function `cos'     incorrect arguments to function `cos'   too few arguments to function `tan'     incorrect arguments to function `tan'   too few arguments to function `asin'    incorrect arguments to function `asin'  too few arguments to function `acos'    incorrect arguments to function `acos'  too few arguments to function `atan'    incorrect arguments to function `atan'  too few arguments to function `ceil'    incorrect arguments to function `ceil'  too few arguments to function `floor'   incorrect arguments to function `floor' incorrect arguments to function `mod'   too few arguments to function `sqrt'    incorrect arguments to function `sqrt'  incorrect arguments to function `pow'   too few arguments to function `min'     incorrect arguments to function `min'   too few arguments to function `max'     incorrect arguments to function `max' abs sin cos tan asin acos atan ceil floor mod sqrt pow min max                           �        incorrect arguments to function `strfind'       incorrect arguments to function `strlen'        incorrect arguments to function `strsub'        incorrect arguments to function `strlower' strfind strlen strsub strlower strupper      Entrada maior que o limite
 Erro ao criar o arquivo "%s"
       Error ao criar o arquivo "%s", atingio o limite de arquivos na entrada de directorio
   Panic: __malloc, sem espaco na tabela de alocacao
      panic: realoc sem espaco, %lx size = %d %d
 PWD BitMAP error
 Not suport BitMAP 4-bit Not suport BitMAP > 8-bit strerrorr
                              (((((�AAAAAABBBBBB                                �Dubug: %s %x %x
        (null)  �o�������h������Di������j�������j������Yk������l������l�������o�������o�������o�������o�������o�������o�������o�������o�������o�������o�������o�������l������vm������(n�������n�������n�������o������.p������.p������.p������.p������p������.p������.p������.p������.p������.p������.p������.p������.p������.p������.p�������o������p������.p������%p������p������.p������p������.p������.p������.p������.p������.p������.p������.p������.p������.p�������o������.p������
p������.p������.p������p������(null) %        :x������gq�������q�������r������Us������t�������t�������t������:x������:x������:x������:x������:x������:x������:x������:x������:x������:x������:x������lu������v�������v������w������w�������x������y������y������y������y�������x������y������y������y������y������y������y������y������y������y������y�������x�������x������y�������x�������x������y�������x������y������y������y������y������y������y������y������y������y�������x������y�������x������y������y�������x������panic: sscanf()
        ��������E����������������������{���������������������������������������������������������������������������������������������������������������������S�����������������������(�������(�������_���������������������������������������z���������������������������������������������������������������������������������������V�������h���������������������������������������h�������������������������������������������������������������������������������_���������������q�����������������������z�������panic: freopen()
 r+ PWD call system funtion error. 
                 $@       �        %lu.%lu                �              �C                                                                        �_�
�@panic: signal()
 panic: sigaction()
 panic: setjmp()  panic: longjmp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �� �   � �   � �     �   � �   �� �    �   � �   X� �   � �   � �   \� �    � �   �# �   �� �   � �   @� �   @ �   (� �   �� �   8� �   H� �   � �     �   `� �                                                   �� �           $� �   h� �   � �   ,� �   �� �           4� �   �� �           <� �   �� �           H� �   �� �           P� �   ~� �           X� �   �� �           `� �   v� �           h� �   �� �           p� �   �� �           |� �   �� �           �� �   �� �           �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   � �   �� �    �   � �   �� �    �   � �   �� �           (� �   �� �           0� �   �� �   @ �   8� �   �� �   p �           �� �           @� �   �� �   � �           �� �           H� �   p� �           P� �   �� �           X� �   �� �           `� �   �� �           h� �   �� �   � �   p� �   �� �                   �� �           x� �   �� �           �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �    � �    �   �� �   �� �    �   �� �   � �    �   � �   �� �           � �   8� �                   &� �                   � �                   � �   @ �   � �   $� �                   �� �   � �    � �   �� �    �   (� �   <� �    �   4� �   �� �    �   <� �   B� �    �   H� �   H� �    �   P� �   �� �    �   X� �   �� �    �   d� �   B� �    �   p� �   $� �    �   x� �   4� �    �   �� �   @� �    �   �� �   <� �    �   �� �   \� �                   Z� �                   J� �                   �� �    �   �� �   h� �                   f� �    �   �� �   R� �    �   �� �   x� �    �   �� �   �� �    �   �� �   p� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �    �   �� �   �� �                   
� �                   |� �                   �� �   P �   �� �   � �    �   �� �   � �    �   �� �   �� �    �   � �   �� �    �   � �   
� �    �   � �   �� �    �   $� �   �� �    �   0� �   � �                   &� �                   �� �    �   <� �   � �    �   H� �   �� �    �   P� �   �� �    �   \� �   �� �           h� �   � �                   � �    �   p� �   8� �                   �� �    �   x� �   �� �           �� �                           �� �   � �   �� �   pU �   pU �                            $ �                           �� �   �� �   �� �   �� �   �� �   �� �   �� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           � �   �f �   �v �   �� �   �� �                           p� �          "{  �   u� �          �{  �   ~� �          �)  �   �� �          d�  �   �� �          |  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  zR x�  ,      @ ���   E�CG����B�A�           L   ����    E�CF���A�(   p   ���Z   E�CG��G�B�A�   $   �   ���l    E�CG��Y�B�A�$   �   "���    E�CG����B�A�$   �   ����    E�CG����B�A�(     l��G   E�CG��4�B�A�   $   @  ����    E�CG����B�A�(   h  ��/   E�CG���B�A�   ,   �  !��   E�CG����B�A�          �  �
��=    E�Ct�      �  ��d    E�CF�T�A�      \��Z    E�CF�J�A�   ,  ���Z    E�CQ�    L  ���J    E�CA� $   l  ����    E�CG����B�A�$   �  ���q    E�CC��b�B�A�$   �  ���    E�CG����B�A�    �  ����    E�CF���A�     U���    E�C��    (  ��@    E�Cw�  8   H  +��C   E�CP�����!�B�B�B�B�A�          �  2��=    E�Ct�     �  O��=    E�Ct�     �  l��0    E�Cg�  (   �  |��   E�CG���B�A�   4     h��M   E�CM�����.�B�B�B�B�A�      H  }��d    E�C[�    h  ���2    E�Ci�      �  ���Z    E�CF�J�A�   �  	��?    E�Cv�  (   �  (��   E�CI�����B�B�A�$   �  ���    E�CG����B�A�$      ����    E�CG����B�A�$   H  ^���    E�CG����B�A�(   p  ! ��o   E�CG��\�B�A�   ,   �  d!��#   E�CL���#�B�B�A�   $   �  PD��|    E�CG��i�B�A�$   �  �D���    E�CG����B�A�$     E��z    E�CG��g�B�A�,   D  lE���   E�CI�����B�B�A�      t  �F���    E�C}�     �  GG��o    E�CE�`�A�   �  �G��_    E�CV� $   �  �G��~    E�CG��k�B�A�      'H��D    E�C{�        KH��D    E�C{�  $   @  oH���    E�CG����B�A�    h  �H��~    E�CF�n�A�$   �  FI���    E�CG��u�B�A�   �  �I��x    E�Co�     �  �I���    E�CF���A�    �  sJ���    E�CF���A�(     K���    E�CI�����B�B�A�    H  �K���    E�CF���A�    l  �L���    E�CF���A�    �  $M���    E�CF���A�$   �  �M���    E�CG����B�A�(   �  {N��   E�CG���B�A�   $   	  mO���    E�CG����B�A�   0	  >P��H    E�C�     P	  fP��H    E�C�     p	  �P��H    E�C�     �	  �P��H    E�C�     �	  �P��H    E�C�     �	  Q��H    E�C�      �	  .Q��|    E�CE�m�A�    
  �Q��p    E�CE�a�A�(   8
  �Q���   E�CG����B�A�   ,   d
  ;T���   E�CI�����B�B�A�   (   �
  �U���   E�CG����B�A�   ,   �
  �X���   E�CI���v�B�B�A�       �
  �Y���    E�CF�v�A�      EZ���    E�CE�}�A�(   8  �Z��a   E�CG��N�B�A�   $   d  �\���    E�CG����B�A�$   �  �]���    E�CG����B�A�(   �  `^��   E�CI�����B�B�A�   �  :_��F    E�C}�  (      `_���   E�CG����B�A�   $   ,  )b���    E�CG����B�A�$   T  �b���    E�CG����B�A�$   |  Wc���    E�CG����B�A�$   �  �c���    E�CC����B�A�$   �  md���    E�CC����B�A�$   �  �d���    E�CC��}�B�A�      He���    E�CE�|�A�$   @  �e��M   E�CE�>�A�      h  �f��v    E�Cm� $   �  *g��5   E�CE�&�A�       �  7h��o    E�CE�`�A�$   �  �h���   E�CE���A�   ,   �  3j���    E�CK������B�B�B�A�   ,  �j��'    E�C^�  $   L  �j���    E�CG����B�A�4   t  �k�� "   E�CM�����"�B�B�B�B�A�   $   �  ����z    E�CC��k�B�A�$   �  ����    E�CG����B�A�$   �  `����    E�CG����B�A�,   $  ώ��F   E�CG��3�B�A�       (   T  ���(   E�CG���B�A�   (   �  ���(   E�CG���B�A�   (   �  ݔ���   E�CJ����B�A�   ,   �  m���p   E�CI���Y�B�B�A�   (     �����   E�CG����B�A�   $   4  F���   E�CG����B�A�(   \  ���'   E�CG���B�A�   (   �  ����   E�CC����B�A�   (   �  ����!   E�CG���B�A�   $   �  ����	   E�CG����B�A�$     m���	   E�CG����B�A�$   0  N���	   E�CG����B�A�$   X  /���	   E�CG����B�A�$   �  ���	   E�CG����B�A�$   �  ���	   E�CG����B�A�$   �  ҫ��	   E�CG����B�A�$   �  ����	   E�CG����B�A�(      ����!   E�CG���B�A�   $   L  ����	   E�CG����B�A�(   t  j���@   E�CG��-�B�A�   (   �  ~����   E�CG����B�A�   (   �  �����   E�CG����B�A�   (   �  r����   E�CC����B�A�   (   $  ���=   E�CG��*�B�A�   $   P   ����    E�CG����B�A�(   x  Ÿ��   E�CG����B�A�   (   �  ����1   E�CG���B�A�   (   �  ����1   E�CG���B�A�   ,   �  ����i   E�CC��Z�B�A�       (   ,  ���Z   E�CG��G�B�A�      X  ���   E�C�   x  ����    E�C��    �  �����    E�C��     �  &���p    E�CF�`�A�$   �  r����    E�CG����B�A�$     1���r    E�CG��_�B�A�(   ,  {���   E�CG��	�B�A�   $   X  k����   E�CF���A�       �  ����    E�CE���A�    �  �����    E�CE���A�   �  ?����    E�C��    �  ����A    E�Cx�        ���i    E�C`�        ,  c���U    E�CL�    L  ����U    E�CL�    l  ����i    E�C`�    �  ���g    E�C^�    �  ]����    E�C�� $   �  $����   E�CE�{�A�      �  ����9    E�Cp�  $     �����    E�CG����B�A�   <  `���^    E�CU� (   \  ����   E�CG���B�A�   (   �  �����   E�CG����B�A�   (   �  %���]   E�CG��J�B�A�   (   �  V���   E�CG��l�B�A�   (     ����D   E�CJ��.�B�A�   (   8  ����:   E�CG��'�B�A�   $   d  ����    E�CG����B�A�   �  �����    E�C��    �  [����    E�C�� (   �  ����   E�CJ����B�A�   (   �  ����i   E�CG��V�B�A�   (   $  ���H   E�CG��5�B�A�   (   P  +���e   E�CJ��O�B�A�      |  d���a    E�CX�    �  ����9    E�Cp�      �  �����    E�CF�w�A�(   �  !���'   E�CG���B�A�   $     ���   E�CE���A�   $   4  �����   E�CF���A�      \  o���    E�C��    |  O����    E�C�� (   �  ���O   E�CG��<�B�A�   $   �  6����    E�CG����B�A�(   �  ����C   E�CG��0�B�A�        ���k    E�Cb� $   <  \����    E�CG����B�A�   d  ����    E�C�� $   �  ����   E�CE��A�   $   �  ����    E�CG����B�A�$   �  ����    E�CG����B�A�(   �  �����   E�CG����B�A�   (   (  #���j   E�CG��W�B�A�       T  a ���    E�CE���� (   x  � ��   E�CG���B�A�       �  ����    E�CE���� (   �  ����   E�CG��q�B�A�   $   �  ���   E�CG����B�A�     ���9    E�Cp�     <  ���+    E�Cb�     \  ����    E�C��     |  L���   E�CE����   �  �
��I    E�C@�     �  ��u    E�CE�f�A�(   �  h���   E�CG����B�A�   (     ���   E�CG����B�A�   $   <  ����    E�CG����B�A�,   d  ���2   E�CG���B�A�          �  ����    E�C��    �  ��w    E�Cn�    �  X��b    E�CY� $   �  ����    E�CG����B�A�$     -��z    E�CG��g�B�A�   D  ��a    E�CX�    d  ����    E�C��    �  :��{    E�Cr� $   �  ���+   E�CF��A�      �  ���6   E�C-�   �  ���L    E�CC� $      ����    E�CG����B�A�   4   z���    E�Cw�    T   ���}    E�Ct� $   t   7��r    E�CF�b�A�    $   �   ����    E�CF���A�       �   ����    E�C��    �   ���3   E�C*�   !  ���7   E�C.�   $!  ���W    E�CN� $   D!  ����    E�CG����B�A�$   l!  Z���    E�CG����B�A�   �!  ����    E�C�� $   �!  t ��V    E�CF�F�A�       �!  � ��P    E�CF�       �!  � ��U    E�CL�    "  !��U    E�CL� $   <"  <!���    E�CG����B�A�$   d"  �!���    E�CG����B�A�$   �"  $"��K    E�CF�{�A�     $   �"  G"��K    E�CF�{�A�     $   �"  j"��S    E�CF�C�A�    $   #  �"���    E�CG����B�A�$   ,#  #��S    E�CF�C�A�    $   T#  0#��K    E�CF�{�A�     ,   |#  S#��[   E�CG��H�B�A�       $   �#  ~$���    E�CG����B�A�$   �#  �$��]    E�CF�M�A�    $   �#  /%��]    E�CF�M�A�    $   $$  d%��K    E�CF�{�A�     $   L$  �%��L    E�CF�|�A�     $   t$  �%��Y    E�CF�I�A�       �$  �%��Y    E�CP� $   �$  &��K    E�CF�{�A�     (   �$  8&���   E�CJ��{�B�A�       %  �.���    E�C��     $   4%  #/���    E�CI���A�       \%  �/��l    E�Cc� (   |%  20���   E�CJ����B�A�       �%  �8���    E�C��     $   �%  a9��   E�CI���A�    $   �%  ::���    E�CI���A�    $   &  �:���    E�CG����B�A�$   D&  �;��\    E�CF�L�A�    $   l&  �;���    E�CG����B�A�$   �&  b<���    E�CI���A�       �&  /=���    E�CI�    $   �&  �=��L    E�CF�|�A�         '  �=��e    E�CF�U�A�    ('  >���    E�CF���A�(   L'  �>���   E�CG����B�A�   (   x'  @��=   E�CG��*�B�A�   $   �'  A��\   E�CE�M�A�      �'  PE���    E�C�� $   �'  �E���    E�CI���A�    $   (  �F���    E�CI���A�       <(  jG���    E�C�� $   \(  �G���    E�CG��z�B�A�   �(  aH��Y    E�CF�       �(  �H��9    E�Cp�  $   �(  �H���    E�CE�q�A�    $   �(  I���    E�CG����B�A�   )  �I��G   E�C>�,   4)  K��u   E�CG��b�B�A�       $   d)  GL��M    E�CF�}�A�     $   �)  lL��O    E�CF��A�     $   �)  �L��L    E�CF�|�A�     $   �)  �L��S    E�CF�C�A�       *  �L���    E�C�    $*  JM���    E�C��    D*  �M���    E�C��    d*  ^N��2   E�C)�$   �*  pQ��U    E�CF�E�A�    $   �*  �Q��U    E�CF�E�A�    4   �*  �Q��L   E�CM�����-�B�B�B�B�A�      +  �S��7    E�C       $   ,+  �S��w    E�CG��d�B�A�(   T+  DT��{    E�CI���d�B�B�A�   �+  �T���    E�C�� $   �+  !U���   E�CE���A�       �+  �W���    E�Cx�     $   �+  HX��\    E�CF�L�A�       ,  |X��5   E�C,�   4,  �[��_    E�CV� ,   T,  �[���   E�CG����B�A�       $   �,  �]��P    E�CF�@�A�    $   �,  �]��Z    E�CF�J�A�    $   �,  �]��^    E�CF�N�A�       �,  ^��4    E�Ck�     -  /^��v   E�Cm�$   <-  �_���    E�CF���A�       d-  `���    E�C�� $   �-  �`���    E�CF���A�       �-  Ra��*    E�Ca�     �-  \a��'    E�C^�     �-  ca��/    E�Cf�     .  ra��;    E�Cr�     ,.  �a��;    E�Cr�     L.  �a��:    E�Cq�     l.  �a��'    E�C^�     �.  �a��9    E�Cp�     �.  �a��9    E�Cp�     �.  �a��<    E�Cs�     �.  b��=    E�Ct�     /  4b��>    E�Cu�     ,/  Rb��n    E�Ce�    L/  �b��;    E�Cr�     l/  �b��9    E�Cp�     �/  �b��9    E�Cp�     �/  �b��9    E�Cp�     �/  c��D    E�C{�     �/  *c��9    E�Cp�     0  Cc��9    E�Cp�     ,0  \c��9    E�Cp�     L0  uc��9    E�Cp�  $   l0  �c��a    E�CF�Q�A�       �0  �c��2    E�Ci�     �0  �c��T    E�CF�   �0  d��X    E�CF�$   �0  Md���    E�CG����B�A�   1  �d��T    E�CF�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    GCC: (Ubuntu 9.3.0-17ubuntu1~20.04) 9.3.0                                        �                  � �                   �                 � �                 � �                  $ �                  T �                    �                	                     ��                     ��_ cole _             ��                )        �           \         �           0    ��                7    ��                >     <"  �   �       C     $#  �   Z      K     ~$  �   l       T     �(  �   /      ^      �� �           c      �� �           h      �� �           m      �� �           r      � �           w      H� �           |    ��                �      T �          �      U �          �     U �          R    U �          �     U �          �     -  �   d       �     h-  �   Z       �     �-  �   Z       �     .  �   J       ^      x� �           c      z� �           h      �� �           m      �� �           r      �� �           w      �� �           �      � �           �      (� �           �    ��                �     PU �          �     XU �          �     �� �          ^      X� �           �    ��                �     `U �          G    x �          �     � �          �     �A  �             �C  �   �           �D  �   �       !    `e �          *    �E  �   o      7    �e �          >    �� �          ^      �� �           c      �� �           h      �� �           m      �� �           r       � �           w      #� �           �      P� �           �      T� �           M     X� �           R     (� �           W     H� �           ]     \� �           c     `� �           i     h� �           o     x� �           u     �� �           {      � �           �     � �           �     � �           �     � �           �     %� �           �     0� �           �     5� �           �   ��                �     $ �    0      �    � �          �    �f �          �    �v �          �    ]�  �   �       �    �  �   a      c     �� �           i     �� �           o     �� �           u     � �           {     *� �           �     A� �           �     P� �           �     x� �           �     �� �           �     �� �           �   ��                �    �� �           [    �# �               �� �               �# �              �� �              �� �          Z    �� �          Y    �� �          K    �� �          J    �� �          ?    �� �          �    �� �              Y�  �   �       %    �  �   �       /    ׏  �   �       :    ��  �   �       E    =�  �   �       T    ܑ  �   �       d    h�  �   �       l    �  �   M      x    @�  �   v       �    ��  �   5      �    �  �   o       �    Z�  �   �      �     � �          �    �� �          �    �� �          �     � �          �    � �          �    � �          �    � �          ^       � �           c      � �           h      (� �           m      ^� �           r      x� �           w      �� �           �      �� �           �      �� �           M     � �           �   ��                �    ļ  �   �       �    `�  �   �       ^       � �           c      (� �           h      L� �           m      U� �           r      ]� �           �   ��                �    =�  �   (          e�  �   (          ��  �   �          I�  �   p      "     � �          .     � �   P       5    ��  �   �      ^      t� �           c      h� �           h      x� �           m      �� �           r      �� �           w      �� �           �      �� �           �      �� �           M     �� �           R     �� �           W     �� �           ]     �� �           c     �� �           i     �� �           o     �� �           u     �� �           {     �� �           �     �� �           �     �� �           �     �� �           �     �� �           �      � �           �     I� �           >     R� �           D     Z� �           J     _� �           P     e� �           V     m� �           \   ��                f    O�  �   !      o    p�  �   	      x    y�  �   	      �    ��  �   	      �    ��  �   	      �    ��  �   	      �    ��  �   	      �    ��  �   	      �    ��  �   	      �    ��  �   !      �    ��  �   	      �    ��  �   @      �    "�  �   �      �    ��  �   �      ^      �� �           c      �� �           h      �� �           m      �� �           r      �� �           w      �� �           �       � �           �      H� �           M     p� �           R     �� �           W     �� �           ]     �� �           c     � �           i     8� �           o     `� �           u     �� �           {     �� �           �     �� �           �      � �           �     (� �           �     P� �           �     x� �           �     �� �           >     �� �           D     �� �           J     � �           P     @� �           V     h� �           �     �� �           �     �� �           �     �� �           �     �� �                �� �           	     �� �                �� �                �� �                �� �           !     �� �           '     �� �           -     �� �           3     �� �           9     �� �           ?   ��                H    �  �   =      Q    T�  �   �       Y    A�  �         a    N�  �   1      k    �  �   1      ^      �� �           c         �           h      P  �           m      y  �           r      �  �           w      �  �           �      �  �           �      �  �           M     �  �           R     �  �           u   ��                |   ��                ^      �  �           c      �  �           h       �           #   ��                �    p� �          ^      p �           c      � �           �   ��                �   ��                ^      � �           �   ��                �   ��                �   ��                �   ��                ^      � �           c      � �           h      � �           �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                   ��                
   ��                   ��                   ��                &   ��                /   ��                8   ��                F   ��                P   ��                Z   ��                d   ��                n   ��                w   ��                �   ��                �    x� �          �   ��                �   ��                �   ��                �   ��                �   ��                ^       �           �   ��                �   ��                �   ��                �   ��                ^      @ �           �   ��                �   ��                �   ��                   ��                   ��                   ��                
   ��                   ��                   ��                "   ��                *   ��                3   ��                <   ��                E   ��                M   ��                T   ��                \   ��                g    �s �   �       ^      X �           ]   ��                j   ��                g    �~ �   �       ^      P �           c      W �           k   ��                v   ��                u   ��                �    �� �          �   ��                   ��                ^   ��                �   ��                ^      P �           �   ��                �   ��                �    ܄ �   e       �    A� �   �       �    � �   �      �    �� �          �    �� �   =      �    �� �          g     � �   �       �   ��                �   ��                �   ��                �   ��                �   ��                ^      X	 �           �   ��                �    �� �   `          ��                ^      j	 �           
   ��                   ��                   ��                "   ��                +   ��                2   ��                >   ��                =   ��                <   ��                D   ��                M   ��                T   ��                [   ��                e   ��                l   ��                ^      m	 �           u   ��                }    �� �          �    �� �          �    �� �   {       �    � �   �       �    Š �   �      �   ��                ^      q	 �           �   ��                ^      �	 �           c      �	 �           h      �	 �           �   ��                �    ɧ �   _       ^      �	 �           c      �	 �           h      �	 �           m      �	 �           �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                   ��                �   ��                   ��                   ��                   ��                #   ��                ^      �	 �           *   ��                0   ��                7   ��                ^      �	 �           >   ��                ^      �	 �           E   ��                ^      �	 �           F   ��                ^      �	 �           8   ��                ^       
 �           ?   ��                ^      
 �           L   ��                ^      
 �           T   ��                ^      
 �           [   ��                ^       
 �           a   ��                j   ��                ^      (
 �           c      9
 �           s   ��                ^      M
 �           c      ^
 �                ��                |    � �           �    ص �   T       �    � �         �    � �   �
      �    �� �   \       �    �< �   �       �    �V �   {       �    .t  �   �       �    �� �          �    �� �   9       �    � �   ;       �    =� �   �       �    �f �          �     O �   �       �    � �   �       
	    �$  �   �       	    �^ �   7      "	    G�  �   �       ,	    �y  �   H           �� �   �       9	    �� �          @	    �u �   �      I	    �  �   '      S	    �� �          ^	    �� �   �       e	    � �           m	    n�  �   �      z	    ry  �   H       Q    /8 �   �       �	    � �           �	    �b �   P       �	     j  �   |       �	    t� �   �       �	    +o  �   D       �	      �          �	    ja �   �       �	    �# �          �    � �          �    2� �   �       �	    �� �          �	    �� �          �	    -- �   �      �	    �o  �   �       �	    M� �   U       �	    �,  �   =       
    �H �   u       
    %� �   w       �    ų �   9       #
    �� �   �      *
    J�  �   �      ;
     �          A
    �)  �         �    �� �   9       J
    �� �   ^       R
    � �          \
    �� �          f
    sv  �   �       v
    f.  �   �       �
    �� �   �       �
    �� �   R      �
    �� �          �    ʍ �   �       �
    �f �   [      �
    � �   :      �
    7 �   �       �
    Jz  �   H       �
    �� �           �    �e �   �       �
    �� �          �
    46  �   0       �
    �S �   w       �
    ?E �   �       �
    2L �   �      �
    � �              �� �   L           �� �              �{  �   p       &    O� �   v      
    T� �   �       -    X� �          7    *�  �    "      ?    or  �   �       N    �b �   U       V    8� �   \       ]    |j �   Y       b    �� �   �      h    �5  �   =       u    �� �   M       L	    �i �   K       �     � �          |    � �          �    1�  �   �       �    �E �   �      �    _A  �   Z       �    �� �          �    ˰ �   <       �    � �   �       <	    � �          �    a1  �   �       �    �� �   L      �    � �   G      �    � �          �    � �              s�  �             p �              �  �             �'  �   �       ,    z  �   H       9    � �   ]      P    �8 �   �       Z    �d �   K       a    \� �          p     � �           u    �n  �   ~       �    Nn  �   _       �    �q  �   �       �    �9 �   �      �    PI �   �      �    �� �          �    h �          �    �5  �   =       �       �           �    �p  �   �       �    ^q  �   x       �    �# �          �    �  �   Z          2 �   �           ��  �   A           �Y �   �           �O �   2      !    W�  �   �       )     �  �   '       0    Ƙ �   2      7    :k  �   z       D    � �          I    Ym  �   �       V    "{  �   |       _    �� �   �       f    �z  �   H       v    R�  �   �       ~    !\ �   �       �    m� �   �       �    �� �   O       �    �� �   5      �    *�  �   i       �    � �   P       �    ׄ  �   �           [t �   �       �    �  �   �       �    MU �   z       �    G  �   #      �     �   �      �    � �          m     ` �           �    72  �   @       �    |c �   �           �� �              �� �   �          #j �   Y           E' �   9       &    � �   �      /    � �          5    (� �   �      }    S� �   9       :    � �          @    @� �          I    �� �          P    J�  �   z       ~     T �           U     �          [       �           b     � �          k     ` �           q    2` �   �       x    ~ �   9       �    ��  �   g       t    ֲ �   D       �    �� �          �    ,� �   '       �    D� �   >       �    �� �   T       �    @� �   �      �    �# �          �    ,b �   V       �    �Z �   �       �    ��  �   U       �    7 �         �    �� �   n       �    2[ �   }       �    �6 �   �       �    �T �   �           Y� �   9             �              �� �   S           O; �   j      "    15 �   k       -    :
 �              T �           9    �� �          ?    �%  �   �       N    �u  �   �       ]    �_ �   W       d    �t  �   �       u    7  �   H      �    #S �   �       �    � �   �       �    �5 �   �       �    7 �          �    �. �          �    C  �   �       �    ` �          �    � �   X       �    ��  �   �       �     �   �       �    �h �   ]       �    @ �          �    � �   D      �    �~  �   �      	     �               � �   �          �  �   �      #     U �   )       �    �` �   �       +    �k  �   �      4    �&  �   G      C     � �   p      K    d �   �       �     � �           Q    B� �   9       ^    Xp  �   ~       m    �� �   ;       w    0T �   b       ~    (� �          �    J�  �   �       �    ��  �   F      �    �j �   K       �    � �   *       �    �0  �   �       �    �d �   K       �    \� �   �       q    S� �   /       �    9�  �   r       �     � �           �    0� �          �    {� �   �       �    �� �          �    �� �   a       �    ,+ �         8    Je �   S       �    E �   +       �    w2  �   C          ��  �   �          �  �   F           9�  �   �           Fu �   l       �    ��  �         $    (V �   �       +    ��  �   i      7    7s  �   �       �    � �   9       F    ��  �   �      _    �H �   I       e    �� �          j    " �   e      v    �@  �   d       }     T �           �    +� �   9       �    �f �   K       A	    1 �         �    u= �         �    c� �   Z       �    �/  �   �       �    hX �   6      �    |  �   �      �    �� �   9       �    Ŭ �   �       �    _� �   2       �    �� �   �       �    � �          �    8� �          �    � �   i      �    �f �          �    c/  �   q           �\ �   �       
    `� �   �           ��  �   �           �� �               ( �   '      �    r� �   �       �     � �           )     � �   �       1    @� �          7    5f �   S       =    ��  �   p       D    @� �   @      H    N   �           V    ��  �   �      a    �2 �   C      m    �� �   :       v    :� �   u      |    ~�  �         �    � �   �       �    /i �   ]       �    H� �          �    |9  �   M      l     ` �           �    Ĉ �   \      �    �i �   L       �    � �   Y       [       �           �    �� �   �      �    �/ �   �       �    � �   7       �    �� �   �      �    P� �          �    � �          �    oo  �   D       �    �& �   a       �    �� �   U           -A  �   2       �
    �C �             [w  �             ~' �   �       �    P? �   �      $    =�  �   i       .    �� �   ;       5    q] �   3      <    `   �   �      A    �> �   �       R    �Y �   L       Y       �           `    'c �   U       h    �D �   9       l    d6  �         r      �   �           2� �   '       Z       �           �    � �   ^       �    � �   �       k    � �   4       �    �U �   a       �    .h �   �       �    d� �   9       �    �j  �   �       �      �   �       �    =W �   +      �    �A  �   ?       �    �z  �   H       �    `� �          �    � �   =       �    d�  �   �      �    � �          �    �m  �   o            k �   �          �[ �   r           ��  �   U       *    K� �   L       /    yx  �   �       @    �0 �   O      H    3�  �   �        lib/setup.asm HEADER_MAGIC HEADER_FLAGS header crt0.c hash.c head present freelist firstnode .LC0 .LC1 .LC2 .LC3 .LC4 .LC5 inout.c nfuncstack fp usererror fileinput fileunput stringinput stringunput .LC6 .LC7 lex_yy.c ncform_sccsid opcode.c base lua_strconc lua_tonumber lua_convtonumber cvt.1965 lua_tostring s.1970 startcode.2115 .LC8 .LC9 .LC10 .LC11 .LC12 .LC13 .LC14 .LC15 .LC16 .LC17 .LC18 .LC19 .LC20 .LC21 .LC22 table.c tablebuffer constantbuffer stringbuffer arraybuffer lua_marktable lua_pack y_tab.c mainbuffer maincode basepc code_byte code_word code_float incr_ntemp incr_nlocalvar incr_nvarbuffer align_n code_number lua_localname lua_pushvar lua_codeadjust lua_codestore msg.2023 yyv yys yypv yyps yystate yytmp lua.c callfunc execstr iolib.c io_readfrom io_writeto io_read buildformat buffer.1817 f.1818 io_write .LC23 .LC24 .LC25 .LC26 .LC27 mathlib.c math_abs math_sin math_cos math_tan math_asin math_acos math_atan math_ceil math_floor math_mod math_sqrt math_pow math_min math_max .LC28 .LC29 .LC30 .LC31 .LC32 .LC33 .LC34 .LC35 .LC36 .LC37 .LC38 .LC39 .LC40 .LC41 strlib.c str_find str_len str_sub str_lower str_upper file.c cfs.c alloc_spin_lock pipe.c path.c gui.c font8x16.c window.c bmp.c font.c border.c memcmp.c memcpy.c memset.c strcasecmp.c strcat.c strchr.c strcmp.c strcpy.c strcspn.c string.c strlen.c strncasecmp.c strncmp.c strncpy.c strpbrk.c strrchr.c strsep.c strspn.c strtok.c last.1481 strstr.c strdup.c memmove.c strcoll.c strerror.c ctype.c tolower.c toupper.c stdio.c fopen.c fclose.c fflush.c fputc.c fgetc.c fgets.c fputs.c fread.c fwrite.c remove.c rewind.c fseek.c feof.c ftell.c vfprintf.c vf vsprintf.c vsnprintf.c sn_buf putchar.c sscanf.c perror.c vfscanf.c character _buf.1638 fvalue _buf.1650 ungetc.c getchar.c freopen.c tmpnam.c _tmpnam rename.c itoa.c i2hex.c malloc.c calloc.c free.c realloc.c lldiv.c strtol.c atoi.c atol.c strtoul.c exit.c getenv.c qsort.c qscmp qses qsexc qstexc qs1 system.c strtod.c ftoa.c _precision atof.c strtof.c strtold.c abs.c ltoa.c utoa.c srand.c errno.c gmtime.c localtime.c strftime.c clock.c math.c pow.c sqrt.c atan.c acos.c asin.c floor.c ceil.c exp.c locale.c signal.c setjmp.c _GLOBAL_OFFSET_TABLE_ longjmp read_directory_blk yysvec drawstring strcpy lua_pushcfunction yyprevious log setjmp lua_nstring clean_blk_enter lua_hashcreate strtok_r lua_parse lua_isnumber stdout vsprintf io_remove lua_ntable ungetc pwd_ptr mathlib_open lua_isnil argv strerror lua_markstack utoa_r lua_getcfunction __m_i memmove lua_string yymorfg __tm __realloc_r lua_getfield atol lua_errorfunction __window_puts getenv yyexca lua_findconstant errno lua_next strtold yyerrflag _infinity lua_storeglobal lua_openfile qsort yycrank yyfnd fgets file_update file_read_block lua_istable yytext yyolsp lua_lasttext memcpy __window_clear BitMAP2 lua_table perror yytchar lua_obj2number ltoa_r lua_debug yyparse lua_pushnumber tolower system feof yyact lua_setunput malloc fs_directory lua_createarray __window_putchar yyoutput lua_nconstant ldexp vsnprintf lua_pushfunction strtoul itoa __pipe__ lua_nfile stdgetc_r yysptr lua_addfile lua_hashmark lua_isstring update_directory_entry _drawline fflush lua_linenumber argc lua_copystring lua_getstring lua_pushnil drawrect BitMAP yylineno yybgin lua_setinput eh_frame lua_getglobal lua_pop lua_constant stdputc_r upath tell_r strncasecmp border write_r yywrap strtol lua_dostring user lua_getparam lua_type rename lua_iscfunction flush_r strrchr utoa calloc strtod rewind_r atof lua_markobject seek_r strcat lua_execute read_directory_entry yynerrs lua_popfunction debug_o yyout yychk fseek __free_block_r open_dir yyval ftoa stdin font8x16 yyleng test __m_c _start obj_list __end strstr write_blk get_file_name yylstate atan2 signal yyr1 lua_array strcoll strncmp write_sector draw_char_transparent strncpy put_pixel strcasecmp log10 _BLK_ realloc drawchar path_count open_file_r yylsp lua_hashdelete lua_pushobject strtok lua_pushuserdata remove_blk memcmp sscanf getfilename file_close pipe_write lua_strdup yytop sigaction read_r file_write_block fread _ctype open_file lua_findsymbol addr yyr2 search_blk_null yyextra lua_call lua_hashdefine yyvstop fopen sysgettmpnam lua_getindexed localtime memset pwd lua_createstring main ftell srand lua_error fclose getchar close_r __data ptr_mouse2 yyestate __free_r update_window lua_reportbug lua_filename getkeyw _vsputs_r strcmp strlib_open lua_pushstring lua_findenclosedconstant color yyin remove_file yyback __bss fgetc drawchar_trans strtof lua_openstring strcspn lua_print ltoa setlocale yydebug stderr create_file lua_narray lua_closefile strsep yypgo getkey yysbuf __malloc_r yymatch mouse fputc open_r A__ call_function iolib_open getpathname strftime i2hex io_execute lldiv fwrite __window yylook vfscanf rewind freopen yydef pipe_read exit yypact pipe_r yylval lua_getuserdata __block_r atoi yyinput lua_storefield __heap_r assert_fn gmtime strspn ctr0 drawstring_trans strlen __code toupper wcl yylex filename_cmp clock read_super_block strchr fputs lua_dofile lua_file strchrnul yyunput lua_isuserdata lua_debugline frexp lua_nextvar yychar lua_getnumber vfprintf strpbrk read_sector free lua_storeindexed setpath yyerror  .symtab .strtab .shstrtab .text .data .got .got.plt .data.rel.local .data.rel .bss .eh_frame .comment                                                                                  �           �                            !              � �    �      P                              '               �         �                              ,             � �   �                                  5             � �   �                                   E              $ �    $      0                              O              T �    T      �                             T                �    `      @                             ^      0                �     *                                                   0�     K         �                	                      H�     P                                                   ��     g                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ELF          >       �   @       8�         @ 8  @  
                 �      �                                      �      �   x        0	                   P      P
 �    P
 �    0       0             Q�td                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��  ���_ cole _          �      �            �
 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           I��H�pF
 �   L�H�PF
 �   H�H�   �   L�H�  �   L�#H�  �   L�+�   �����H��H��H��H��L�������UH��AWSH��@��H�����I��     L�H�}�H�u�H�U�H�M�L�E�L�M�H���������H�H�U�H�H�	     H�E�H�H�E�H��	     H�H��	     H�H� H��H� 	     H�H��	     H�H��H��	     H�H��	     H�H�@H��H��	     H�H�E�H��	     H�H�E�H��	     H�H�E�H��	     H�H�	     H�H��H��	     H�I�߸    H�O������H���H��	     H�    H���������H�H� H��H��	     H�H���������H�H� H��H���������H�H� H�։�I��H���������H��ЉE�E��I��H�r�������H��АH��@[A_]���UH��AWAUATSH��0��H�����I�     Lۉ}�H�u��}�9H�E�H� H��H� �������H�<I�߸    H�~�������H��Ҹ   �  H�E�H��H� H�F�������H�4H��I��H���������H���H�E�H�}� u/H�P�������H�<I�߸    H�~�������H��Ҹ   �  H�Eغ   �    H��I��H���������H���H�E�H��I��H�Y�������H��ЉEԋEԉ�I��H�3�������H���H�E�H�Eغ    �    H��I��H���������H��ЋU�H�M�H�EȾ   H��I��H�V�������H��ЉE�H�E�H��I��H�8�������H���H�X������H��ЋU�H�Eȉ�H��H��������H��Ѕ�t/H�p�������H�<I�߸    H�~�������H��Ҹ   �  �}�~
H�E�H�@�2H��������H��Ѕ�tH���������H��H���������H�H���������H�4H��I��H���������H���H�E�H�}� u/H���������H�<I�߸    H�~�������H��Ҹ   ��   H��������H���A��H�Z������H���A��H��������H��Ѕ�t�   ��   H�E�E��D��H���������H�43H��I�߸    I�ߛ������I�A��H�K������H���A��H��������H���H��H�E�H��D��   I��H���������H���H�E�H��I��H�8�������H���H��������H��и    H��0[A\A]A_]���UH��H����H�����I��     L؉}��}� x�}��   �E���������    ����UH��H��8��H�����I�?     L�H�}�H�E�H��� ���E�H�Eȋ@�E��E�E�H�UȋR�U�E�H�UȋR�U�E�H�UȋR�U�E�H�UȋR�U�E�H�UȋR�U�E��uhH�EȋH�E�H�����H�U�H��� �H�E�H����H�U�H��� �H�E�H����H�U�H��� �H�E�H�����H�Eȉ��  H�Eȋ ���耉E��U��E��i�5  �E܋E�i��  �E�ЉE��E�iв����E�ЉE�U�E��i�h	  �E܋E�i������E�ЉE�E�i�O����E�ЉE�U��E�ЉE܋E�)E��U�E��i�T  �E��E�i�8����E�ЉE��E�i�   �E�ЉE�U��E�ЉE��E�)E��U�E�ЉE�E�)E�U܋E�ЉE�E�)E܋U��E�ЉE�E�)E��U��E��i��   �����E��E�+E�i��   �����E��U�E������H�Eȉ�U�E��H�E�H������U��E��H�E�H������U܋E��H�E�H������E�+E��H�E�H������E�+E���H�E�H������E�+E���H�E�H������E�+E���H�E�H���������UH��SH��H��H�����I�x     L�H�}�H�u��U�H�E�H�耋 ���E�H�E����   �E�E�E�H�U��R@�U�E�H�U��R �U�E�H�U����   �U�E�H�U����   �U�E�H�U��R`�U�E؅�uSH�E�� �� ���耉�H�l�������H������E��E�   ��E���H�E���E�H�HE��m��}� u��  H�E�� ��    �E�U�E��i�5  ���EԋE�i��  �E�����E�E�iв����E�����E��U܋E��i�h	  ���EԋE�i������E�����E܋E�i�O����E�����E؋U�E�ЉEԋE�)E�U�E��i�T  ���E��E�i�8����E�����E�E�i�   �E�����E�U�E�ЉE��E�)E�U��E�ЉE܋E�)E��UԋE�ЉE؋E�)EԋU�E�ЉE�E�)E�U�E��i��   �����E�E�+E�i��   �����E�U؋E�����耉�H�l�������H���H�U���E�H�HE��U�E�����耉�H�l�������H���H�U���E�H�HE��U�E�����耉�H�l�������H���H�U���E�H�HE��UԋE�����耉�H�l�������H���H�U���E�H�HE��E�+E����耉�H�l�������H���H�U���E�H�HE��E�+E����耉�H�l�������H���H�U���E�H�HE��E�+E����耉�H�l�������H���H�U���E�H�HE��E�+E����耉�H�l�������H���H�U��H��H[]���UH��H����H�����I��     L؉}�}� �<  �    �  H�        �T��TH�        ��� ���р��H�        ��� H�        ��� �JH�        ��� ��  H�        H�TH�JH�        H�L0��U�H�        �T�J�H�        �LH�        ��� �JH�        ��� H�        ��� �����U�	�H�        ��� �}���)  H�        �T���  H�        H�TH�JH�        H�L0��U�H�        �T�J�H�        �L�U����   ��   ���   '����   ���   uH�        �D    �   �U����   ���   tH�        �   �hH�        ��� �����U�	�H�        ��� H�        ��� �JH�        ��� ���H�        �   H�        ��� 9U������H�        ��� H�        ��� +E�����E�   �������!�����UH��SH����H�����I�     Lۉ}�H�        ��� 9E�~�E��H� �������H���H�        ��� +E�H�        ��� �H��[]���UH��SH����H�����I��     Lۉ}�E��H� �������H��ЉE�E��H���������H��ЋE�H��[]���UH����H�����I�4     L�H�        ��� �с��   H�        ��� �]���UH��H����H�����I��     L؉}�H�        H�L�U�Hc�H�H�        H�LH�        �T+U�H�        �TH�        �T+U�H�        �TH�        �T��yH�        �   �����UH��H����H�����I�1     L�H�}�H�E�� ������H�E�H��� ��	�����UH��S��H�����I��     L�H�        �D��H�        �   �{H�        H�DH��H���������H�����H�        �DH�        �TH�        �D9�~H�        �   ��   H��������H���[]���UH��S��H�����I�&     L�H��������H���H�        �D��H��������H��А[]���UH��AWSH�� ��H�����I��     L��E�    �E�    H��������H���H�        �D��H�        �   �  H�        H�D� <tH�        �   �f  H�        H�DH��H��H���������H�����H�        �DH�        H�DH��H��H���������H�����H�        �DH�        H�DH��� ��H�        �D0�   H��������H���H�        �D0��t��tH�        �   �  �H�        �LH�        �T0����9�}H�        �   �Q  �E�    H�X       H�H�E���  H�        H�D� ��H�E؉H�        H�DH��� ����H�E؉PH�E؋@��uH�        �   ��  H�E؋PH�E؋@��!Ѕ�tH�        �   �  H�        H�DH��� ������H�E؉PH�E؋@��uH�        �   �a  H�E؋PH�E؋@��!Ѕ�tH�        �   �4  H�        H�DH��� ��H�E؉PH�E؋@%�   ��tH�        �   ��  �   H��������H���H�        ���   H�E؋@�   �����	�H�        ���   H�E؋@9E�}
H�E؋@�E�H�E؋@9E�}
H�E؋@�E�E�H�E�0H�        �D09E��$���H�        �D0��u7H�X       H�H�E��E�   �E�E�H�E؋U�PH�E؋PH�E؉P�E��    H�        �T(�E��    H�        �T,H�        �TH�        �D(Ѓ�H�        �t(�����H�        �T H�        �TH�        �D,Ѓ�H�        �L,�����H�        �T$�E�    H�X       H�H�E��m  H�        �TH�E؋@�ЋE�Ѓ���}��H�E؉PH�E؋@��%�����H�E؉PH�        �TH�E؋@�ЋE�Ѓ���}��H�E؉PH�        �T H�        �D(��H�E؋@��}��H�E؉PH�E؋@��H�E؋@9E�uH�E؋@��"H�E؋@9E�tH�        �   �M  H�E؋HH�        �T$H�        �D,��H�E؋@��}�����I��H�3�������H���H�U�H�B(H�E�H�@(H��uH�        �   ��   �E�H�E�0H�        �D09E��|���H�        �D0����   H�        �TH�        �D��H�        �D0��I��H�3�������H���H�        H��� H�        H��� H��uH�        �   � H�        �D��H��������H���H�� [A_]���UH��ATSH��0��H�����I��     L�H��������H����"  H�        H�D� ���E��E�%�   ��tH�        �   �#  �E�����tH�        �   �  �E���E����E��E�   �7H�        H�T�E�H�HЋU�r��H�     Hc�Hو�E��}�~ÿ   H��������H��ЋE�H�H��H���  H�        H�H�H�E��E�   �E�E��E�   ��   �}�E��H�     H�H�����Ẽ}� ��   H�        �D9E�~H�        �   �  �   +E�Ủ����)E�}� yH�        �   ��   �E�    �IH�        H�T�E�H�H�D� �E�E���E��H�EЈH�E�D�`H�E��m��}� uރE��E�;E�|��Ẻ�H��������H������E��}�������H�E��  H�E��E�P��U��u�H�        �D�������H�        �D��tH�        �   �H��0[A\]���UH��SH����H�����I�"     L�H��������H�����   H�        H�D� ���E�E�%�   ��tH�        �   ��   H�        ���   �E��   �����	�H�        ���   �E�H�H��H���   H�        H�H�H�E��E�    �2H�        H�D�U�Hc�H��HЋU�Hc�H�U�H�� ��E��}�?~ȿA   H��������H���H�        �D��@����H�        �D��tH�        �   �H��[]���UH��S��H�����I��     L�H��������H���H�        �D��H�        �   �VH�        H�DH��H���������H�����H�        ��� H�        �D��H��������H���[]���UH��SH�� ��H�����I�     L�H�}�H�uؿ   H� �������H��ЉE�E�H�H� H�E�H�� ���E��}� uH�        �   �    �   �E���H���������H��ЋE�H�H� H�E�H��@���E�H�}� t�E��H�E؈�E���E��}� u�    �E�E���H�e�������H��ЉE�E����   �����9E�}�E���������Ѓ�E�E�H�� []���UH��AWSH�� ��H�����I��      L�H�}�H�u��E� �E�    �   �    H��     H�<I��H��{������H���H�E؋@ H�H��H���  H�        H�Hо    H��H���������H���H�U؋R$�H�E؉P$H�E؋P$H�E؋@H�        H�H�H��H�H�   � ����H�        ��� H�E؋@H�H��H���  H�        H�H�H�E�H��H��H���������H��ЉE��E����   �E�������u�E�<�tH�        �   �b  �E�������E�}�?~H�        �   �6  H�E؋PH�        �E�H�Hc�H�H��H�H�H�   � ��H� ��������U�Hc�H�����E�H�        Hc�H��t  H��H�H�H����}�>��������E�    �?�E�H�Ht  H��    H�        H�H�H��H��H���������H��ЃE��}�?~��E�    �XH�E؋@�U�Hc�H�U�H�4�U�Hc�H��t  H��    H�        H�H�H�J��H��H�{�������H��ЃE��}�~�H�� [A_]���UH��SH��8��H�����I��      L�H�        ��� �E��E�    H��������H���H�        �DH�        �T0���9�}H�        �   ��  H�        H�D� ��H�        �D09�tH�        �   ��  �   H��������H����E�    H�X       H�H�E���   H�        H�D� ��H�Eȋ 9�tH�        �   �X  H�        H�DH��� ��%�   ��tH�        �   �   H�        H�DH��� ����H�EȉP H�        H�DH��� ��������H�EȉP�   H��������H��ЃE�H�E�0H�        �D09E�����H�        H�D� ��u4H�        H�DH��� <?uH�        H�DH��� ��tH�        �   �@  H�        �D��H��������H����E�    �E�E��E�    H�X       H�H�E��   �E�    �   �E�    �qH�E�H�P(H�Eȋ@�E���E��H�Eȋ@��H�Eȋ@�E���E����H�H�H�E�H��H��H��������H���H�        ����r  �E�H�Eȋ@9E�|��E�H�Eȋ@9E��f����E�H�E�0H�        �D09E��:����E�H�        �D 9E�|"�E�    �E�H�        �D$9E���   H�        ��� ��������m��}� �����H���������H��п   H�e�������H��ЉE�E�%��  =��  u�E��9E�tH�        �   �z�Eԃ����E�H�        ��� �E��E�    �1H�        �E�Hc�H��H�H�H��H�H�H��\�     �E��}�~������H�        �   ��H��8[]���UH��AWATSH��H��H�����I���      L�H�}�H�E��@���E�H�E��PH�E��@�����I��H�3�������H���H�E�H�}� uH�        �   �  H�E�H�@(H�E�H�E�H�E�H�E��@�E��  H�E�� ��iЋ   H�E�H��� ��k��Ѓ�@����H�l�������H���H�UЈH�E�� ��k�hH�E�H��� �Љ��Ѝ�    ЍH�E�H��� ������)���Ѓ�@��H�U�L�b��H�l�������H���A�$H�E�� ��k�H�E�H��� ��k�m�H�E�H��� �Љ������ȃ�@��H�U�L�b��H�l�������H���A�$�E�    �J  �E�Hc�H�E�H�� �Љ�����؋U�Hc�H�JH�U�H����k�oE�H�H�HH�E�H�� ��k�E�H�H�HH�E�H�� ������)���Ѓ�@���U��Hc�H�JH�U�L�$��H�l�������H���A�$�E�Hc�H�E�H�� ������)E�H�H�HH�E�H�� ��k�E�H�H�HH�E�H�� ��k�o��E�H�H�PH�E�H�� �Љ������ȃ�@���U��Hc�H�JH�U�L�$��H�l�������H���A�$�E��E�;E������H�E��@H�HE�H�E��@�H�HE�H�E�H��� ��k�H�E�H��� ��k�m�H�E�H��� �Љ������ȃ�@��H�U�L�b���H�l�������H���A�$H�E�H��� ��k�hH�E�H��� �Љ��Ѝ�    ЍH�E�H��� ������)���Ѓ�@��H�U�L�b���H�l�������H���A�$H�E�H��� ��iЋ   H�E�H��� ��k��Ѓ�@��H�U�L�b���H�l�������H���A�$�m��}� �P���H�E��@� H�E��PH�E��PH�E��PH�E�H�@(H��I��H�Ͻ������H���H�E�H�U�H�P(H��H[A\A_]���UH��AWSH��@��H�����I���      L�H�}�H�E��@�E�H�E��@�EЋE���E�H�E��PH�E��@�����I��H�3�������H���H�E�H�}� uH�        �   �9  �E�    ��  H�E�H�P(�E�H�H�H�E�E�Hc�H�E�H�H�E�H�E�� ��iЋ   �E�Hc�H�E�H�� ��k��Ѓ�@����H�l�������H���H�U���E�H�HE�H�E�� ��k�h�E�Hc�H�E�H�� �Љ��Ѝ�    ���E�Hc�H�E�H�� ������)�ȃ�@����H�l�������H���H�U���E�H�HE�H�E�� ��k��E�Hc�H�E�H�� ��k�m��E�Hc�H�E�H�� �Љ������ȃ�@����H�l�������H���H�U���E�H�HE��E�H�HE�H�E��@���E��!  �E���Hc�H�E�H�� �Љ������H�U����k�o��E�Hc�H�E�H�� ��k���E�Hc�H�E�H�� ������)�ȃ�@����H�l�������H���H�U���E�H�HE��E���Hc�H�E�H�� ������)�H�E�� ��k���E�Hc�H�E�H�� ��k�o��E�Hc�H�E�H�� �Љ������ȃ�@����H�l�������H���H�U���E�H�HE��E�H�HE�m��}� ������E�H�HE�H�E�� ��k��E���Hc�H�E�H�� ��k�m��E���Hc�H�E�H�� �Љ������ȃ�@����H�l�������H���H�U���E�H�HE�H�E�� ��k�h�E���Hc�H�E�H�� �Љ��Ѝ�    ���E���Hc�H�E�H�� ������)�ȃ�@����H�l�������H���H�U���E�H�HE�H�E�� ��iЋ   �E���Hc�H�E�H�� ��k��Ѓ�@����H�l�������H���H�U���E��E�;E�����H�E��@� H�E��PH�E��PH�E��PH�E�H�@(H��I��H�Ͻ������H���H�E�H�U�H�P(H��@[A_]���UH��AWAVAUATSH��X��H�����I��      L��E�    H�X       H�H�E��  H�E��PH�        �D9�}H�E�H��H�o������H���H�        �����  H�E��PH�        �D9�}H�E�H��H�������H���H�        �����  H�E��PH�        �D9��Y���H�E��PH�        �D9��<���H�E��PH�        �D9�|H�E��PH�        �D9�}H�        �   �
  �E�H�E�0H�        �D09E��^���H�        �D0����  H�        H��� H�E�H�        H�D`H�E�H�        H���   H�E�H�        H���   H�E�H�        �D�E��O  �E�    ��   �E�Hc�H�E�H�� ����A�ċE�Hc�H�E�H�� ��D�p��E�Hc�H�E�H�� ��D�x�Ai�g  D�����L�m�I�UH�U���H�l�������H���A�E AkƨA�Ai�I���Ѓ���L�m�I�UH�U���H�l�������H���A�E Ai��  D�����L�e�I�T$H�U���H�l�������H���A�$�E�H�        �D9E�� ���H�        �DLH�HE�H�        �D|H�HE�H�        ���   H�HE��m��}� ������
  H�        �TDH�        �DL9���   H�        H�T`H�        �DLH�H�H�E�H�        H�T`H�        �DDH�H�H�E�H�        �DH���E��\H�        �DD��H�M�H�E�H��H��I��H�={������H���H�        �DLH�HE�H�        �DDH�HE��m��}� u�H�        �DDH�        �DL����H��X[A\A]A^A_]���UH��AWH����H�����I���      Lغ� �    H�        H�<I��H��{������H��ѐH��A_]���UH��AWSH����H�����I�@�      L��E�    �rH�        �E�Hc�H��H�H�H��H�H�H��`H� H��t?H�        �E�Hc�H��H�H�H��H�H�H��`H� H��I��H�Ͻ������H��ЃE��}�~�H�        H��� H��t'H�        H��� H��I��H�Ͻ������H���H�X������H��АH��[A_]���UH��SH����H�����I�B�      L�H�}�u�H��������H���H�        H�E�H�D�E�%�����H�        �TH�        �D��
�   �  H�        H�D� �Љ�H�        H�DH��� ���	Є�t
�   ��  �   H��������H����\  H�        �D��~H�        H�D� <�t
�   �  �   H��������H���H�        H�DH��� ��=�   ;=�   ��   -�   ����   ��H��    H� �  H�H��  H�>��=�   tb�rH�&�������H����   H�/�������H����   H���������H����tH�4�������H����bH��������H����PH���������H����>H�        H�DH��� ��%�   =�   uH���������H�����   �iH�        ��������H�        ���tH�        ��3H�        �    �    H��������H���H�        �H��[]���UH����H�����I���      L�H�        �D]���UH����H�����I�n�      L�H�        �D]���UH����H�����I�>�      L�H�        �D0������]���UH����H�����I��      L�H�        �T0��uH�        H�D`�H�        H��� ]���UH����H�����I���      L�H�        �LH�        �T��H�        �D0��]���UH��AWSH����H�����I�T�      Lۉ}�H�u�H�E�� ��H�E��@9�sH�E��P#H�E��@9�r"H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@��u)H���������H�H��E�H�։�H��������H���H�E�H�PH�E��@#��H�H�E�H�PH�E�H�@�U�H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  H�E��@��u0H���������H�H� H��t�E�����I��H�Pm������H��ЋE�H��[A_]���UH��H����H�����I���      L�H�}��E�    H�E�@��u]H�E�@'�PH�E�P'��H�E�P#H�E�@'9�r�H�E�H�PH�E�@'��H��H�H�E�H�PH�E�H�@� ���E��   H�E�@��tH�E�@��uiH�E�@#��u������ZH�E�P'H�E�@#9�r������AH�E�H�PH�E�@'��H�H�E�H�PH�E�H�@� ���E�H�E�@'�PH�E�P'�E�����UH��H����H�����I���      L�H���������H�H� H�E��E�    H�E��@��uWH�E��P#H�E��@'9�w�    �AH�E�H�PH�E��@'��H�H�E�H�PH�E�H�@� ���E�H�E��@'�PH�E��P'�E�����UH��H����H�����I�7�      L�H���������H�H� H�E��E�    H�E��@��uXH�E��@'�PH�E��P'��H�E��P#H�E��@'9�r�H�E�H�PH�E��@'��H��H�H�E�H�PH�E�H�@� ���E��E�����UH��AWH��(��H�����I���      L�H�}�H�u�H�U����u�    �(H�M�H�U�H��H��I��H�=5������H���H�E�H�E�H��(A_]���UH��AWSH�� ��H�����I��      L�H�}�H�}� u
������   H�}� tH�E؋@����tH�E��@"<t������zH�E؋@%�   ��u�    �cH�E؋@#H�U؋J�    ��E�H�E؋@��@��u�U�H�E؉�H��I��H��?������H���H�E�H��I��H��<������H��ЉE�E�H�� [A_]���UH��AWSH����H�����I�4�      L�H�}�H�}� u������0H�E�H��H��������H���H�E�H��I��H��=������H���H��[A_]���UH��AWSH�� ��H�����I���      Lۉ}�H�u�H�}� u
�������  H�EЋ@��u
�    �  H�EЋ@��tH�EЋ@��tH�EЋ@��u!H�UЋE�H�։�H��������H����y  H�EЋ@����unH�EЋP#H�EЋ�+  9�wYH�EЋ�+  ��tKH�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��E�U�H�EЉ�H��I��H��>������H����H�EЋ@����H�EЉPH�EЋ@#H�UЋJ�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U܈H�E�� ��H�EЋ@��9�r3H�EЋ@����H�EЉPH�E�f�   H�E�H��H��������H���H�EЋ@#�PH�EЉP#H�EЋP#H�EЋ�+  9�vH�EЋ�+  �PH�EЉ�+  H�EЋ@���H�EЉP�    H�� [A_]���UH��AWH��(��H�����I���      L�H�}�H�}� u
������  H�E؋@��u
�    �v  H�E؋@��tH�E؋@��tH�E؋@��u"H�E�H��H��������H��ЉE�E��0  H�E؋P#H�E؋�+  9�r
������  H�E؋@����ulH�E؋P#H�E؋�+  9�wWH�E؋�+  ��tIH�E؋@����H�E؉PH�E؋@#H�U؋r�    ���E�U�H�E؉�H��I��H��>������H���H�E؋@#H�U؋J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@� ���E�H�E�� ��H�E؋@��9�rH�E؋@����H�E؉PH�E�f�   H�E؋@#�PH�E؉P#�E�H��(A_]���UH��SH��H��H�����I���      L�H�}ȉuĉU�H�M�H�}� u�    �y�E�    H�E�H�E��E�    �FH�E�H��H�K!������H��ЉE؃}��u�E�    �u��4H�E�H�PH�U��U؈�E��E��E��E��E�9�w��E�    �u�H��H[]���UH��SH��H��H�����I��      L�H�}ȉuĉU�H�M�H�}� u�    �l�E�    H�E�H�E��E�    �9H�E�H�PH�U�� ���E�H�U��E�H�։�H�/������H��ЃE��E��E��E��E�9�w��E�    �u�H��H[]���UH��H����H�����I�e�      L�H�}�H�u��U�}�tZ�}�|�}� t�}�t�nH�E���H�E��P#H�E���H�E��P'�RH�E��@#H�U��H�E��P#H�E��@'H�U��H�E��P'�(H�E���+  H�U�)Љ�H�E��P#H�E��P#H�E��P'�H�E��@#H�U��J�    ��Љ�H�E�f��    ����UH��H����H�����I���      L�H�}�H�}� u�    �	H�E��@#������UH��H����H�����I�F�      L�H�}�H�}� t7H�E��@'    H�E��P'H�E��P#H�E�f�   H�E��@����H�E��P������UH��H��(��H�����I���      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H��(��H�����I���      L؉}�u�H�U�H�M��E������   �E�H�u�H�}؉��r�E��E�����UH��H����H�����I�3�      L�H�}��E�_   �(�E�Hc�H�E�H�� < u�E�Hc�H�E�H��  �m��}� y����    ����UH��H����H�����I���      L�H�}�H�E�H�E�H�E�H�E��H�E�� </uH�E�H��H�E�H�E�H�E�� ��u�H�E�����UH��H��0  ��H�����I�`�      L�H������H������H������H�E�H������H�E�H������H�E��E�    �?H�E�� ��u�E�Hc�H�E�H��  �H�E�H�PH�U��U�Hc�H�U�H�� ��E��}�_~��E�    �-H�E�H�PH�U��H�E�H�PH�U�� 8�t�   ��E��}�_~͸    ����UH��SH�� ��H�����I�{�      L�H�}�H�u�H�E؋PH�E؋@ЉE�E�H�U����H�@	     H�H�¾   H�&������H��ЉE�}� t
�������   �E�    ��   �E�%�  ��H�@	     ��H؋���uf�E�%�  ��H�@	     ��H��������E�H�U����H�@	     H�H�¾   H�l&������H��ЉE�}� t������r�E��m�E�%�  =�  uE�E��E�H�U����H�@	     H�H�¾   H�&������H��ЉE�}� t�������E�H�E؋@$9E����������H�� []���UH��H����H�����I���      L؉}��u�H�U�H�M�    ����UH��AWSH��0��H�����I���      Lۉ}�H�u�H�U�H�EȋPH�Eȋ@ЉE�H�Eȋ@ �E܉E�ЉE�   �    H�@	     H�<I��H��{������H����E�    �B�U�E�Љ�H�EЋ ��H�@	     H��   H�l&������H��ЉE��}� u�E�H�EȋP �E�9�w���H��0[A_]���UH��H����H�����I���      L�H�}�H�u�H�U��R��H�U����H�U�H��H��   I�&������J� ������UH��AWSH��`��H�����I�o�      L�H�}�H�u�H�U�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H�3�������H���H�E�H�E�H�E�H�E�H��I��H��\������H��ЉE�H�E��@,�E��9  H�E�H�E��H�E�� </uH�E��  H�E��H�E�H�E�� ��u׋U�H�E��@ H�M��	��H�M���H�&������H��ЉE؃}� t#H�E�H��I��H�Ͻ������H��и    ��   �E�    �f�E���Hc�H�E�H�H�E�H�E��@a��t5H�E��@b����@��t#H�E�H�U�H��H��H��'������H��ЉE���E������}� t�E��}�?~����}� u+�}�?%H�EЋ@k�E�H�E��@ �E؉E�ЉE�m��	�E�    �
�}� �����H�E�H��I��H�Ͻ������H��ЋE�H��`[A_]���UH��AWSH��P��H�����I�Z�      L�H�}�H�u�H�U��M�L�E�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE�    I��H�3�������H���H�E�H�Eغ    �    H��I��H��{������H��ЋU�H�E��@ H�M��	��H�M؉�H�&������H��ЉE�}� t#H�E�H��I��H�Ͻ������H��и������   �E�    �T�E���Hc�H�E�H�H�E�H�E��@a��t#H�E�H�U�H��H��H��'������H��ЉE���E������}� t�E��}�?~����}� u:�}�?4�E���Hc�H�E�H�H�EȺ�   H��H��I��H�={������H�����E�����H�E�H��I��H�Ͻ������H��ЋE�H��P[A_]���UH��AWSH��P��H�����I���      L�H�}�H�u�H�U�H�E���C  ��u
������	  H�E���C  ��@v/H�0�������H�<I�߸    H�~�������H��Ҹ������  H�E��PH�E��@ЉE�H�E���?  H�E��@ �ЋE�ЉE�    I��H�3�������H���H�E�H�Eغ    �    H��I��H��{������H��ЋU�H�E��@ H�M��	��H�M؉�H�&������H��ЉEԃ}� t!H�E�H��I��H�Ͻ������H��ЋE��  H�E���C  ��H��H��H�E�H�H�E�H�EȺ`   �    H��I��H��{������H���H�E�H��+H��H�*'������H���H��H�E�H��H��I��H�F~������H����E�    �"H�UȋE�H����uH�UȋE�H�� �E��}�_~�H�E��@` H�E���+  H�EȉPo�U�H�E��@ H�M��	��H�M؉�H�l&������H��ЉE�H�E�H��I��H�Ͻ������H��ЋE�H��P[A_]���UH��AWSH��`��H�����I�3�      L�H�}�H�u�H�U��S  I��H�3�������H���H�E�H�EкS  �    H��I��H��{������H���H�E��PH�E��@ ��H�EЉP�    I��H�3�������H���H�U�H�BH�E��PoH�EЉ�+  H�E��PH�EЉ�/  H�E��P H�EЉ�3  H�E��H�EЉ�G  �    I��H�3�������H���H�U�H��K  H�E�H��K  �    �    H��I��H��{������H���H�E��@k�E�    I��H�3�������H���H�E��E������E�    �E�    ��  �   I��H�3�������H���H�U�H��K  �M�Hc�H��H�H�H�E�H��K  �U�Hc�H��H�H� H�E�H�E��   �    H��I��H��{������H����E�    �<  H�E��@ �E��H�E��@�H�E��P�E�H�H�4�    H�E�H�ʉH�EЋ�;  �PH�EЉ�;  �E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E�;E�ts�E�H�U����H�U�H��H�¾   H�&������H��ЉE��}� t:H�E�H��I��H�Ͻ������H���H�E�H��H��=������H��и    �   �E��E�H�E��@�����E�    ��U�E�H��    H�E�HЋ �E�}��u	�E�������E��}��  ������}��t�E��}��  � �����H�E�H��I��H�Ͻ������H���H�E�H��`[A_]���UH��AWSH��p  ��H�����I���      L�H������H�������   I��H�3�������H���H�E�H�E�H�E�H�E�H   H�E�H������H�E�H��H��I��H�rZ������H���H�U�H�E�H��H��I��H� ]������H��п�   I��H�3�������H���H� 	     H�H� 	     H���   �    H��I��H��{������H��п   I��H�3�������H���H�E�H�EȺ   �    H��I��H��{������H���H�E�H�E�H�E��   �    H��I��H��{������H����E�    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ����    Hǅ ���    Hǅ���    Hǅ���    Hǅ���    Hǅ ���    Hǅ(���    Hǅ0���    Hǅ8���    Hǅ@���    HǅH���    HǅP���    HǅX���    Hǅ`���    Hǅh���    Hǅp���    Hǅx���    H�E�    H�E�    H������H������H��H��I��H�F~������H���������<wt������<au�E�   H�E��@   H�E��     H�U�H�E�H��H��H�$+������H��ЉE�}� t_H� 	     H�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H��и    �  H�E�H�U�H�M�H�E�H��H��H��+������H��ЉE��}� u_H� 	     H�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H��и    �  H�EȋU��P,H� 	     H�H�M�H�U�H�u�I�ȹ    H��H��-������H��ЉE�}����   �}� tqH� 	     H�H������H�U�H�u�A�    H��H�RD������H���H� 	     H�H������H�U�H�u�I�ȹ    H��H��-������H��ЉE�}� ��   H� 	     H�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H��и    ��  �}� t_H�E�H��I��H�Ͻ������H���H� 	     H�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H��и    �r  H� 	     H�H�U�H�M�H��H��H��1������H���H�E�H�}� ��   H� 	     H�H��H�E�H��+�`   H��H��I��H�={������H���H�E�H��+H��H��&������H���������<wt������<+t������<au
H�E��@"�H�E��@"H�E��@   H�EȋP,H�E���?  H� 	     H��PsH�E���C  ������<auH� 	     H��PoH�E��P#H�E�H��I��H�Ͻ������H���H� 	     H�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H���H�E�H��p  [A_]���UH��AWSH��@��H�����I�p�      L�H�}��   I��H�3�������H���H�E�H�E�   �    H��I��H��{������H���H�E�H�E�H�E�   �    H��I��H��{������H���H�E��@   H�E��     H�U�H�E�H��H��H�$+������H��ЉE܃}� t H�E�H��I��H�Ͻ������H��и�����AH�U�H�M�H�E�H��H��H�a/������H��ЉE�H�E�H��I��H�Ͻ������H��ЋE�H��@[A_]���UH��AWSH�� ��H�����I�6�      L�H�}�H�E�H�@H��I��H�Ͻ������H����E�    �TH�E�H��K  �U�Hc�H��H�H� H��t?H�E�H��K  �U�Hc�H��H�H� H��I��H�Ͻ������H��ЃE��}��  ~���H�E�H��K  H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H���H�E�    �    H�� [A_]���UH��H�� ��L�����I�9�      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H�&������I� ������UH��H�� ��L�����I�e�      M�H�}�u�H�E苐;  �E�9�vH�}� u
������   H�E�H��K  �E䍈�  ��H���
H�H��H�H� H�E��E����%�  )�H�H��    H�E�HЋ �E�H�E�H�H�U�H�E苀3  H�u苶G  ����H�l&������I� ������UH��AWSH��   ��H�����I���      L�H��x���H��p�����l����   I��H�3�������H���H�E�H�E�H�E�H�E�H   H�E�H��x���H�E�H��H��I��H�rZ������H���H�U�H�E�H��H��I��H� ]������H��п   I��H�3�������H���H�E�H�EȺ   �    H��I��H��{������H���H�E�H�E�H�E��   �    H��I��H��{������H���H�E��@   H�E��     H�U�H�E�H��H��H�$+������H��ЉE��}� t_H� 	     H�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H��и�����-  H�E�H�U�H�M�H�E�H��H��H��+������H��ЉE��}� u_H� 	     H�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H��и�����  H�EȋU��P,H�EȋPH�Eȋ@ЉE�H�EȋP,H�Eȋ@ �ЋE�ЉE��    I��H�3�������H���H�E�H�E��    �    H��I��H��{������H��ЋU�H�Eȋ@ H�M��	��H�M���H�&������H��ЉE��E�    �E�    �   �E���Hc�H�E�H�H�E��E�;�l���}~H�E��@a��ta�E���Hc�H��p���H�H�E���   H��H��I��H�={������H��ЋE���Hc�H��p���H�H��H��&������H��ЃE����E��}�?�e�����H�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H��ЋE�H�Đ   [A_]���UH��AWSH��`��H�����I���      L�H�}�H�u�H�U�H�M�D�E�H�E�H�E�H�Eغ�   �    H��I��H��{������H���H�E�H��H�*'������H���H��H�E�H��H��I��H�F~������H����E�    �"H�U؋E�H����uH�U؋E�H�� �E��}�_~�H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉEп    I��H�3�������H���H�E�H�EȺ    �    H��I��H��{������H��ЋU�H�E��@ H�M��	��H�Mȉ�H�&������H��ЉEă}� t!H�E�H��I��H�Ͻ������H��ЋE���  �E�    �$�E���Hc�H�E�H�H�E�H�E��@a��t�E��}�?~���H�E��@a���G  �}�?�=  �U�H�E؉PsH�E��@a��E���H�E؈PbH�U�H�E�H��H��H�x(������H���H�U؉BkH�E؋@k���uOH�E�H��H�L�������H�<I�߸    H�~�������H���H�E�H��I��H�Ͻ������H��и   ��   �E���@��t$H�E؋@kH�U�H�M�H�Ή�H�;*������H���H�M�H�E຀   H��H��I��H�={������H��ЋU�H�E��@ H�M��	��H�Mȉ�H�l&������H��ЉEĐH�E�H��I��H�Ͻ������H��и    �JH�E�H��I��H�Ͻ������H���H�E�H��H�p�������H�<I�߸    H�~�������H��Ҹ����H��`[A_]���UH��AWSH��P��H�����I�6�      Lۉ}�H�u�H�U��    I��H�3�������H���H�E��E�    �E��E��E������E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��E��E܋E�;E���   �}� tV�E�H�U����H�U�H��H�¾   H�l&������H��ЉẼ}� t#H�E�H��I��H�Ͻ������H��и�����?  �E�H�U����H�U�H��H�¾   H�&������H��ЉẼ}� t#H�E�H��I��H�Ͻ������H��и������   �E��E�E��E��E�   H�E��@�����E�    ��U�E�EȋE�H��    H�E�HЋ �E�E�H��    H�E�H��     �}��uL�E�H�U����H�U�H��H�¾   H�l&������H��ЉE̐H�E�H��I��H�Ͻ������H��ЋE��6�E��    H�E��p�Ⱥ    ����H�E��@�H�E��@ЉE��Y���H��P[A_]���UH��AWSH��   ��H�����I��      L�H��h����   I��H�3�������H���H�E�H�E�H�E�H�E�H   H�E�H��h���H�E�H��H��I��H�rZ������H���H�U�H�E�H��H��I��H� ]������H��п   I��H�3�������H���H�E�H�E��   �    H��I��H��{������H���H��p���H�E�H�E��   �    H��I��H��{������H���H�E��@   H�E��     H�U�H�E�H��H��H�$+������H��ЉE�}� t<H�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H��и    ��  H�E�H�U�H�M�H�E�H��H��H��+������H��ЉE��}� u<H�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H��и�����d  H�E��U��P,H�E��PH�E��@ЉE�H�E��P,H�E��@ �ЋE�ЉE��    I��H�3�������H���H�E�H�E��    �    H��I��H��{������H��ЋU�H�E��@ H�M��	��H�M���H�&������H��ЉE�}� tSH�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H��ЋE��l  �E�    �   �E������E���Hc�H�E�H�H�E�H�E��@a��t!H�E�H�U�H��H��H��'������H��ЉE�}� u9H�E��@a �U�H�E��@ H�M��	��H�M���H�l&������H��ЉE�}� ��E��}�?�k����}� tPH�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H��ЋE��uH�E��@kH�U�H�M�H�Ή�H��G������H��ЉE�H�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H���H�E�H��I��H�Ͻ������H��ЋE�H�Đ   [A_]���UH��H����H�5����I���      Lމ}�E�E��}� u�E��   �E����rH�P	     H�H�P	     H�����UH��H����H�����I�+�      L�H�}��   H�E�H���r�����UH��AWH����H�����I��      L�H�@	     H�H�U�H�H	     H�    H�      �    H�M�   �    H��I��H��{������H��ѐH��A_]���UH��AWSH��P��H�����I�h�      Lۉ}��u��}� u
�    ��  H�H	     H�H=�   v%H���������H�<I�߸    H�~�������H��ҐH�      ���u�H�      ��PH�      ��E����E�E�%�  ��t�E��E�    �E�    �E�    �}� t�E��   �E�   �K  �}��  �=  H�@	     H�H�E�H�E�    �E�    �  H�E؋@����   H�E؋@9E���   H�E�H�H�E؋@��H�H�E�H�E؋@+E���H�E؉PH�E؋P�E��H�E؉PH�E�H�E�H�@	     H�H�E��E�    �mH�E؋@��tH�E��E��WH�E�H�E�H�E�H�E�H�E�H�@H�PH�E�H�PH�E��@   H�E�H�U�H�H�E��U��PH�E�H�U�H�P�E���!�}��   ~��H�E��E��}��   ������E�   ���}� ��   H�@	     H�H�E��E�    �~H�E؋@��tH�E��E��hH�E�H�E��E��H�hN������H���H�E�H�E�H�U�H��E��E���H�E��PH�E��U��P�E���+E���H�E��PH�E�H�@   ��}��   �u���H�      �    H�H	     H�H�PH�H	     H�H�E�H��P[A_]���UH��SH��(��H�����I�C�      L�H�}�H�}� ��  �H�      ���u�H�      ��PH�      �H�E�H�E�H�@	     H�H�E��E�    �M  H�E�H� H9E�tH�E��E��2  H�E�H�E�H�H	     H�H�P�H�H	     H�H�E؋@��uH�E�H��H��N������H����   H�E؋@��uH�E�H�@H�E�H�E�H�@H�P�H�E�H�PH�E�H�@H��tH�E؋@����   H�E�H�@H��uRH�E�H� H��H��N������H���H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    H�E�H�     H�E��@    H�E��@    H�E��@    H�E�H�@    ��}��   �������H�      �    ��H��([]���UH��AWH��H��L�����I�A�      M�H�}��u�H�E�    �E�    H�}� u�E��   ��H��O������I� ���8  �H�      A� ��u�H�      A� �PH�      A� H�@	     I� H�E�H�E�H�E��E�    �   H�E�H� H9E�t
H�E��   H�E�H�E��E�   H�E��P�E��=   v@H�H	     I� �U�H�E�H��H� �������I�< M�Ǹ    I�~�������M�A����H�E�H� H�E�H�E��P�E��H�E��P�E��}��   �X���H�      A�     �}� u�E��   ��H��O������I� ���H�E�H��HA_]���UH��H�� ��H�����I���      L�H�}�H�u��E�    H�E�H�E��   H�E�� ��H�E��@9�sH�E��P#H�E��@9�rH�E��@#    H�E�f�   H�E�H�PH�E��@#��H�H�E�H�PH�E�H�PH�U�H�U�H�R� �H�E��@#�PH�E��P#H�E��P#H�E���+  9�vH�E���+  �PH�E���+  �E��}��E����E�����UH��H�� ��H�����I���      L�H�}�H�u��E�    H�E�H�E�H�E��@'�PH�E��P'H�E��P'H�E��@9�rH�E��@'   �H�E��P#H�E��@'9�r�H�E��@'�P�H�E��P'�JH�E�H�PH�E��@'��H�H�E�H�PH�E�H�PH�E�H�HH�M���H�E��@'�PH�E��P'�E��}�~��E�����UH��AWSH��0��H�����I���      L�H�}�H���������H�H� H�E�H�E�H�E�H�E�H��I��H�"�������H��ЉE�H�E�H��I��H�"�������H��ЉE؋U܋E��=   ~
������   H�E�� </uH�E��E�H�HE�H�m�H�E�� </tH�E�H�E�H�PH�U�� /�H�E�H�U�H�E�H��H��I��H�F~������H���H�E�H��I��H�"�������H��Љ�HE�H�m�H�E�� </u	H�E��  �H�E�H�E��  �    H��0[A_]���UH��AWSH����H�����I�k�      L�H���������H�H� H��I��H�"�������H��Ѓ�w
�    �   H���������H�H� H�E�H�E�H��I��H�"�������H��Љ�HE��H�E�H�P�H�U��  H�E�� </u�H���������H�H� H��I��H�"�������H��Ѓ�vH�E��  �    H��[A_]���UH��AWSH��0��H�����I��      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
�    ��  H�E�H��I��H�"�������H��ЉE�E�H�H�P�H�E�H�� </u�E�H�H�P�H�E�H��  �}� 
�    �  �}���   H�E�H��� <:u%H�U�H�E�H��H��I��H�F~������H����K  H�,�������H�<I��H���������H���H��H�E�H��H��I��H�F~������H���H�E�H��I��H�"�������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H�F~������H����   H�,�������H�<I��H���������H���H��H�E�H��H��I��H�F~������H���H�E�H��I��H�"�������H��ЉE�H�E�� </t�E�Hc�H�E�H�� /�E��E�Hc�H�E�H�H�E�H��H��I��H�F~������H���H�E�H��0[A_]���UH��H����H�����I�?�      L�H�}�H�E�H�E�H�}� u�    �+�E�    �H�E�� </u�E�H�E�H�E�� ��u�E�����UH��AWSH��0��H�����I�Ѣ      L�H�}�H�u�H�E�H�E�H�E�H�E�H�}� tH�}� u
������   H�E�H��I��H�"�������H��ЉE�E�H�HE�H�m��H�E�� </tH�m�H�E�� ��t�E�P��U�����H�E�H�U�H�E�H��H��I��H�F~������H���H�E��  �    H��0[A_]���UH��H��0��H�����I��      L�H�}�H�u��U܉M�L�E�H���������H�H� H�E��E�H9E�}?H�E��@��H9E�}0H�E�H�E��E�H�E�H��H�E�H�H��    H�E�HE؉������UH��SH��@��H�����I�U�      Lۉ}ԉuЉỦM�L�E�L�M�f�E�  H�E�H�@H�E�H�E��@�E�}�u�E�    �E�    �   f�E� H�E��@�EȉE��H�H� H�E�H�� f�E�H�E�� ���E��J�E�f#E�f��t5�UЋE��Hc��UԋE��H�H�}��M�U�I��H��H�^������H���f�e�m��}� y��E�H�E��@9E��b�����H��@[]���UH��AWSH��0��H�����I�>�      Lۉ}܉u؉UԉM�D�E�L�M��E�    �X�E�    �CH�E�L��   �M�H�E��P�u؋E��Hc��}܋E��H�H��I��H�^������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I���      Lۉ}܉u؉UԉM�D�E�L�M��E�    �p�E�    �[H�E�H��   �E��E�i��E��A��H�E��P�M؋E��Hc��M܋E��H�I��D��H��I��H�^������H��ЃE��E�;E�|��E��E�;E�|���H��0[A_]���UH��AWSH��0��H�����I�Ȟ      Lۉ}܉u؉UԉM�D�E�L�M��}� �[  �}� �Q  �E�    �>H�E�L��   �M�H�E��P�E�Hc��}܋E��H�H��I��H�^������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E����Hc��}܋E��H�H��I��H�^������H��ЃE��E�;E�|��E�    �AH�E�H��   �M�H�E��P�u؋E��Hc��E�H�I��H��I��H�^������H��ЃE��E�;E�|��E�    �FH�E�L��   �M�H�E��P�u؋E��Hc��}܋E����H�H��I��H�^������H��ЃE��E�;E�|���H��0[A_]���UH��AWSH��@��H�����I��      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}��  �E�    ��   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��   �E�f#E�f��tDH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�^������H����BH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�^������H���f�e�m��}� �[����E�H�E��@9E��	�����H��@[A_]���UH��SH��8��H�����I���      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H��b������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I���      Lۉ��uȉUĉM�D�E�L�M�f�E�f�E�  H�E�H�@H�E�f�}���   �E�    �   f�E� �U�H�E��@�ЋE��H�H� H�E�H�� f�E�H�E�� ���E��W�E�f#E�f��tBH�EH��   H�E�P�MċE��Hc��MȋE��H��M�I��H��I��H�^������H���f�e�m��}� y��E�H�E��@9E��T�����H��@[A_]���UH��SH��8��H�����I�ۙ      L�H�}؉uԉUЉM�D�E�L�M��E�    H�E�H�E��^H�E���E�P�U��ȉʋEԍ4H�E�H�PH�U�� f���L�E��}ȋM̋U�H���uM��A����H��d������H���H��H�E�� ��u���H�]�����UH��AWSH��@��H�����I��      L�H�}ȉuĉU��M�D�E�D�M�H���������H�H� H�E�H�E�H   � �? �    H��I��H��{������H����E�    �U�H�E��P4�UH�E��P8�UH�E��P<H�E��@H   H�E��@L   H�E��P<H�E��PP�UH�E��PTH���������H�H��H�E�H�PXH�E��@D    H�E��PDH�E��P@�U�H�E��P�U�H�E��P�U�H�E��P �U�H�E��P�U H�E��P`�} u�E�   H�E��@�P�H�E��P(H�E��P�E�)ЍP�H�E��P$H�E��@0   �E����H�E��P,H�E��@��H�E��@��H�E�I���Ѻ    �    I��H�uw������H���H�E��@4��H�E��@����H�E�I��A�ȹ   �   �   H��_������H��Ѓ}� u:H�E��@����H�E�I��A���� �   �   �   H��_������H����8H�E��@����H�E�I��A���� �   �   �   H��_������H��Ѓ}� t}H�E��@����H�U��E�I��A���� ����   �   H��_������H���H�E��@4��H�E��@���ƋE��H�U�I��A�ȹ   ��ƿ   H��_������H���H�E��@8A��H�E��@$��H�E��@(��H�E��@,��H�E��@0��H�E�I��H��_������H���H�E�H��I��H�"�������H������E�H�E�H�pHH�E��@��E܉������)Љ�H�E�H���u�I��A���� ������   ��H��H�f������H���H��H�E��@����H�E�I��A�    �   �   �   H�)a������H���H�E�H�PHH�E��@��H���u�I��A���� ������   �ƿX   H��d������H���H��H�E�H�PHH�E��@��(H���u�I��A���� ������   �ƿ-   H��d������H���H��H�E�H�e�[A_]���UH��AWSH��0��H�����I���      L�H�}�H�u�H�E��P0H�E��@Ѓ�P�E�H�E��P,H�E��@Ѓ��E��E�P   �E�   �E�    �E���� H�E�H��I��H�"�������H��ЉE�H�E�L�@H�M؋U܋E���������p��E�<�E��������ƋE���)ƋE��H�E�H���u�M��A�ȉщ�H��H�=d������H���H���H�e�[A_]���UH��H����H�����I���      L�H�}��   H�E�H���r�����UH��H����H�����I�\�      L�H�}������UH��H����H�����I�1�      L�H�}�H�U��BD    H�U��JDH�U��J@H�U��R8A��H�U��R$��H�U��R(A��H�U��R,��H�U��R0��H�U�I��D��I��_������J��А����UH��SH��(��L�����I���      Mډ�f�E�H���������I�H� H�E�H���������I�H��H�E�H�PXH�E�@(�P�H�E�@H���к    ��E�H�E�@$�P�H�E�@L���к    ��E�H�E�P<H�E�PPH�E�PD�E�9�rH�E��@D    H�E�@@�PH�E�P@H�E�P@�E�9�r9H�E��@D    H�E�PDH�E�P@H�E�H��H��l������I����E��  f�}���   H�E�@D����   H�E�@D�P�H�E�PDH�E�H�xHH�E�pTH�E�@PH�U�J,H�U�RLA��H�U�R@A��ʃ���H�U�J0H�U�RHA��H�U�RDA��ʃ�A��H���u�I��A������D�޿    H��b������I���H����   f�}�	uH�E�@D�PH�E�PD��   f�}�
u!H�E��@D    H�E�@@�PH�E�P@�   f�}���   H�E�H�xHH�E�pTH�E�PPH�E�H,H�E�@LA��H�E�@@A��ȃ���H�E�H0H�E�@HA��H�E�@DA��ȃ�A���E�H���u�I��A���щ�D�މ�H��b������I���H��H�E�@D�PH�E�PD�E�H�]�����UH��H����H�����I�ޏ      L؉}�H���������H�H� H�E��U�H�E��P<�����UH��SH��(��H�����I���      L�H�}�H�}� t=H�E�H�E��&H�E�H�PH�U�� f�����H�Pm������H���H�E�� ��u���H��([]���UH��AWSH��P��H�����I��      L�H�}��u��U��M�L�E�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H�0�������H�<I�߸    H�~�������H��Ҹ�����6  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H�>�������H�<I�߸    H�~�������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�V�������H�<I�߸    H�~�������H��Ҹ   ��   �E�    �   �E�    �   �}� tNH�E�H��   H�E��P�M��E���E��Hc��M��E���E��H��M�I��H��I��H�^������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�^������H��ЃE��}� �U����E��}� �;����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��P��H�����I�;�      L�H�}��u��U��M�D�E�L�M�H�E�H�E�H�E�H��6H�E�H�EЋ@
��H�E�H�H�E��E�    H�E�� f=BMt/H�0�������H�<I�߸    H�~�������H��Ҹ�����3  H�EЋ@�E��  �E�    ��  H�E��@f��wtH�E��@f��u/H�>�������H�<I�߸    H�~�������H��Ҹ   ��  �E��P�U�Hc�H�E�H�� ��H��    H�E�HЋ %��� �E��   H�E��@f����   H�E��@f��u%�E��P�U�����Hc�H�E�HЋ %��� �E��ZH�E��@f�� u�E��P�U���Hc�H�E�HЋ �E��/H�V�������H�<I�߸    H�~�������H��Ҹ   ��   �E�    �   �E�    �   �}� tKH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�^������H����IH�E�L��   �M�H�E��P�u��E�ƋE��Hc��}��E�ǋE��H�H��I��H�^������H��ЃE��}� �X����E��}� �>����E�H�EЋP�E�9�������m��}� ������    H��P[A_]���UH��AWSH��0��H�����I�X�      Lۉ}܉u؉U�H�M��E�    �   �E�    �t�U�������E��H���������H�Hڋ��E�}� tBH�E�H��   H�EȋP�MԋE��Hc��M؋E��H��M�I��H��I��H�^������H��ЃE��}�~��E��}��o�����H��0[A_]���UH��AWSH��@��H�����I�|�      Lۉ}̉uȉUĉM�L�E��E���� �E�``` �E���� �EĉE��ẺE܋E��E؋EȉEԋE؍P��E��xH�M��E�I��A�    �   ��I��H�)a������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H�)a������H��ЋE؍P��E܍p�E���H�}��M�I��A�ȹ   ��I��H�)a������H��ЋEԍP��E܍pH�M��E�I��A�    �Ѻ   ��I��H�)a������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H�)a������H��ЋEԍP��E܍p�E���H�}��M�I��A�ȉѺ   ��I��H�)a������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H�)a������H��ЋEԍP��E܍p�M��E�ȃ�H�}��M�I��A�ȉѺ   ��I��H�)a������H��ЋEԍP��E܍p�M��E�ȃ�H�M�I��A�    �Ѻ   ��I��H�)a������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H�)a������H��ЋE؍P��M܋E�ȍp��E���H�}��M�I��A�ȹ   ��I��H�)a������H��ЋE؍P��M܋E�ȍp��E���H�M�I��A�    �   ��I��H�)a������H��АH��@[A_]���UH��H��8��H�����I�M�      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �CH�E�H�PH�U�� ���E�H�E�H�PH�U�� ���E�E�+E�E�}� u�}� t
�m��}� u��E�����UH��H��8��H�����I���      L�H�}�H�uЉŰẺE�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M����E��P��U���u�H�E�����UH��H�� ��H�����I�@�      L�H�}���U��E�E��E�H�E�H�E��H�E�H�PH�U��U��m��}� u�H�E�����UH��AWSH��0��H�����I�ۃ      L�H�}�H�u�H�E�H�E�H�E�H�E��E�    H�E�H�PH�U�� ����I��H�V�������H��ЉE�H�E�H�PH�U�� ����I��H�V�������H��ЉEԋE�+EԉE܃}� u�}� t뗋E�H��0[A_]���UH��AWSH����H�����I� �      L�H�}�H�u�H�E�H��I��H�"�������H��Љ�H�E�H�H�E�H��H��I��H�F~������H���H�E�H��[A_]���UH��H�� ��H�����I���      L�H�}�u�H�E�H�E��H�E�� ��9E�uH�E��H�E�H�E�� ��u۸    ����UH��H�� ��H�����I�H�      L�H�}�H�u�H�E�H�E�H�E�H�E��3H�E��H�E�� 8�u!H�E�� ��H�E�� ��Ѕ�u�    �'H�E�H�PH�U��H�E�H�PH�U�� 8�t����������UH��H��0��H�����I���      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E��  H�E�����UH��AWH��(��H�����I�1�      L�H�}؉uԋU��҉Uԃ}� uOH�U�H��I��H�"�������H��҉�H�E�H���   H�E�� ��tH�E�� ��9E�u	H�E��   H�E�H�E؃�H��űE�i��E�H�E�H�E��H�E�H�E� ������H�E� ��!�%������u%H�E� 3E䍐����H�E� 3E���!�%������t�H�E�H�E��H�E�H�E�� ��tH�E�� ��9E�u�H�E�H��(A_]���UH��H��@��H�����I��      L�H�}�H�u�H�U�H�U�H�U������   H�U�H�������   H�E�    H�E�    H�E�    H�E�    �H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�t�H�E�H+E��'H�U����H�Uȉ�H��H��~������H���H+E�����UH��H����H�����I��~      L�H�}�H�E�H�E��H�E�H�E�� ��u�H�E�H+E�����UH��AWSH��@��H�����I��~      L�H�}�H�u��U�H�E�H�E�H�E�H�E��E�    �kH�E�H�PH�U�� ����I��H�V�������H��ЉE�H�E�H�PH�U�� ����I��H�V�������H��ЉEԋE�+EԉE܃}� u�}� t
�m��}� u��E�H��@[A_]���UH��H��(��H�����I��}      L�H�}�H�u��U�H�E�H�E�H�E�H�E��}� u)������2H�E�H�PH�U��H�E�H�PH�U�� 8�u�m��}� u����E�����UH��H��8��H�����I�>}      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��E�    �!H�U�H�BH�E�H�E�H�HH�M����E��E�9E�w�H�E��  �E�����UH��AWH����H�����I��|      L�H�}�H�u�H�M�H�U�H��H��I��H��������H��҉�HE�H�E�� ��tH�E���    H��A_]���UH��AWH��(��H�����I�M|      L�H�}؉u�H�U�H��I��H�"�������H��҉E��U�H�E�H�H�E��E�    �H�E�� ��9E�uH�E��H�m��E��E�9E�wڸ    H��(A_]���UH��H��0��H�����I��{      L�H�}�H�u�H�E�H� H�E�H�}� u�    �vH�E�H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u,�}� u
H�E�    �H�E�H���  H�E�H�U�H�H�E���}� u������UH��H��@��H�����I��z      L�H�}�H�u�H�E�H�E�H�E�    H�E�    H�E�    H�E�    H�E�� ��u
�    ��   H�E�H��� ��u+�H�E�H�E��H�E�� 8�t�H�E�H+E��   H�E�H�E�� ��tAH�E�� ���Ћt��H�U���҃��   �������	�T�ЋD�Ѕ�u��H�E�H�E�� ��t/H�E�� �����T��H�E�� �����   �����!Ѕ�u�H�E�H+E�����UH��H��8��H�����I��y      L�H�}�H�u�H�U�H�}� uH�E�H� H�E�H�}� u
�    ��   �H�E�H�PH�U�� ���E�H�E�H�E��
�E�;E�u��H�E�H�PH�U�� ���E��}� uۃ}� uH�E�H�     �    �   H�E�H��H�E�H�E�H�PH�U�� ���E�H�E�H�E�H�E�H�PH�U�� ���E��E�;E�u4�}� u
H�E�    �H�E�H��H�E�H�E��  H�E�H�U�H�H�E���}� u������UH��H����H�����I��x      L�H�}�H�u�H�u�H�M�H�(     H�H��H�(�������H�������UH��AWSH�� ��H�����I�;x      L�H�}�H�u�H�E�H��I��H�"�������H��ЉE��2�U�H�M�H�E�H��H��I��H��z������H��Ѕ�uH�E��H�E�H�E�� ��uø    H�� [A_]���UH��AWSH�� ��H�����I��w      L�H�}�H�E�H��I��H�"�������H��Ѓ��E�E��I��H�3�������H���H�E�H�}� u�    �$�U�H�M�H�E�H��H��I��H�={������H��АH�� [A_]���UH��H��8��H�����I�w      L�H�}�H�uЉU�H�E�H�E�H�E�H�E��U�H�E�H�H�E�H�E�H;E�v[H�E�H;E�sQH�E�H�E��E�HE��H�m�H�m�H�E��H�E��H�E�H;E�u��'H�U�H�BH�E�H�E�H�HH�M���H�E�H;E�u�H�E�����UH��AWH����H�����I�Bv      L�H�}�H�u�H�M�H�U�H��H��I��H��}������H���H��A_]���UH��AWH����H�����I��u      Lډ}�H�p�������H�<I�׸    H�~�������H�������UH��H����H�����I��u      L؉}��U���H���������H�Hc��������t�E� �E�����UH��H����H�����I�Iu      L؉}��U���H���������H�Hc��������t�m� �E�����UH��AWSH��0��H�����I��t      L�H�}ȉuĉU��M��U�H�E�H��H���������H�<I�߸    I�~�������I�A��H�E�H��I��H��������H���H�E�H�E� �E�H�E� 9E�u��H��0[A_]���UH��AWSH�� ��H�����I�Ot      L�H�}�H�u�H�E�� ��u�    �LH�E�� <wuH�E�H��I��H��������H���H�U�H�E�H��H��I��H�f������H���H�E�H�E�H�� [A_]���UH��AWH����H�����I��s      L�H�}�H�U�H��I��H��������H���H��A_]���UH��AWH����H�����I�os      L�H�}�H�U�H��I��H��������H���H��A_]���UH��AWH����H�����I�$s      L؉}�H�u�H�M��U�H�Ή�I��H�/������H���H��A_]���UH��AWSH�� ��H�����I��r      L�H�}�H�}� u������VH�E�H��I��H�K!������H��ЉE�H�E؋@��u+H���������H�H��E�H�։�I��H�/������H��ЋE�H�� [A_]���UH��AWH����H�����I�9r      L؉}�H�u�H�M��U�H�Ή�I��H�Ό������H���H��A_]���UH��AWH����H�����I��q      L�H�}�H�U�H��I��H�!�������H���H��A_]���UH��AWSH��@��H�����I��q      L�H�}ȉu�H�U�H�}� u	H�E��  H�E�H�E�H�E�H�E��E�    H�E�H��I��H�K!������H��ЉEԃ}����   H�E��@��u7�}�u�}� ~+H���������H�H��E�H�։�I��H�/������H��Ѓ}�
tk�E�;E�}E�}�u�}� ~H�E�H;E�vH�m��m��:�}��^���H�E�H�PH�U�UԈ�E��D����}�u�}� ~�m���E��)�������}�~	H�E��  ��Eԉ�H�E�H�E�H��@[A_]���UH��AWSH�� ��H�����I�?p      L�H�}�H�u�H�}� u�    �^�E�    �2�E�Hc�H�E�H�� ��H�U�H�։�I��H�Ό������H��ЃE�H�E�H��I��H�"�������H��ЋU�9�w��E�H�� [A_]���UH��AWH��(��H�����I��o      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I�#������I�A��H��(A_]���UH��AWH��(��H�����I�?o      L�H�}�u�U�H�M�H�M؋U��u�H�}�I��I��#������I�A��H��(A_]���UH��AWH����H�����I��n      L�H�}�H�U�H��I��H�J������H���H��A_]���UH��AWH����H�����I��n      L�H�}�H�U�H��I��H��%������H��ҐH��A_]���UH��AWH��(��H�����I�Kn      L�H�}�H�u��U܋U�H�u�H�M�H��I��H��$������H���H��(A_]���UH��H����H�����I��m      L�H�}�H�}� u������!H�E��P#H�E���+  9�r�������    ����UH��AWH����H�����I��m      L�H�}�H�U�H��I��H�m%������H���H��A_]���UH��AWSH��`  ��H�����I�Jm      L�H������H������H�������E�    �E�    �  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H�5�������H���	E�}���  �E�H��    H�c  H�H�c  H�>��H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E��E�H������H�։�I��H���������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�}� t(H������H�E�H��H��I��H���������H����O  H������H��H���������H�<I��H���������H����   H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �E�H�������E�H�։�I��H�w�������H���H������H������H��H��I��H���������H����w  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������
   H��H��I��H���������H���H������H������H��H��I��H���������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�J� �EċE�H�������   H��H��I��H���������H���H������H������H��H��I��H���������H����  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�EȾ   H��fHn�I��H���������H���H������H������H��H��I��H���������H����]  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eк
   H��H��I��H�I�������H���H������H������H��H��I��H���������H����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ
   H��H��I��H���������H���H������H������H��H��I��H���������H�����  H������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H������H�Eغ   H��H��I��H���������H���H������H������H��H��I��H���������H����G  H�������@=�   w3H������H�PH�������@��H�H�������R�JH�������J�H������H�@H�HH������H�J� �E�H������H�E�   H��fHn�I��H���������H���H������H������H��H��I��H���������H����   H������H�ƿ%   I��H���������H��ЋE�Hc�H������H�� ��H������H�։�I��H���������H����4�E�Hc�H������H�� ��H������H�։�I��H���������H��ЃE��E�Hc�H������H�� ��������    H��`  [A_]���UH��H����H�����I��d      L؉��E��E�    �E��S��%wa��H��    H��[  H�H��[  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I�d      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��H�� ��H�����I�*c      L�H�}�H�u�H�E�H�E�H�E�H�E��H�U�H�BH�E�H�E�H�HH�M���H�E�� ��u�H�E�����UH��AWSH��  ��H�����I��b      L�H������H������H��x����E�    H������H�E�f�E�  �E� �E�    �/  �E�    �E�Hc�H������H�� ������%��  �E��E�Hc�H������H�� ������lu�E��E�   �E�Hc�H������H�� ����H��������H���	E܃}���  �E�H��    H�fZ  H�H�[Z  H�>��H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E��E�H�U�H�E�H��H��H�ʜ������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H�}� t'H�U�H�E�H��H��H�ʜ������H���H�E��e  H�E�H���������H�4H��H�ʜ������H���H�E��7  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E�H�������E�H�։�I��H�w�������H���H������H�E�H��H��H�ʜ������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������
   H��H��I��H���������H���H������H�E�H��H��H�ʜ������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�J� �E��E�H�������   H��H��I��H���������H���H������H�E�H��H��H�ʜ������H���H�E��3  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�E��   H��fHn�I��H���������H���H������H�E�H��H��H�ʜ������H���H�E��x  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�E��
   H��H��I��H�I�������H���H������H�E�H��H��H�ʜ������H���H�E���  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ
   H��H��I��H���������H���H������H�E�H��H��H�ʜ������H���H�E��  H��x���� ��/w0H��x���H�PH��x���� ��H�H��x�����JH��x����
�H��x���H�@H�HH��x���H�JH� H�E�H������H�EȺ   H��H��I��H���������H���H������H�E�H��H��H�ʜ������H���H�E��e  H��x����@=�   w3H��x���H�PH��x����@��H�H��x����R�JH��x����J�H��x���H�@H�HH��x���H�J� �E�H������H�Eо   H��fHn�I��H���������H���H������H�E�H��H��H�ʜ������H���H�E��   H�E�H���������H�4H��H�ʜ������H���H�E�fǅ����  �E�Hc�H������H�� ������H������H�E�H��H��H�ʜ������H���H�E��8�E�Hc�H������H�� �E�H�U�H�E�H��H��H�ʜ������H���H�E��E��E�Hc�H������H�� �������H�E��  H�U�H������H)�H��H�Ā  [A_]���UH��H����H�����I��Y      L؉��E��E�    �E��S��%wa��H��    H�S  H�H��R  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I�:Y      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H�6�������L��Љ�<�����<���Hc�H�����H��  ��<���H���   A_]���UH��AWH���   ��L�����I�9X      M�H����������H�����H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H����������H�����H��M��H���������L��Љ�<�����<���H���   A_]���UH��AWSH��0��H�����I�NW      L�H�}؉u�H�U�H�M��}�   v
�    �   H�U�H�E�H��H�@     H�<I��H�6�������H��ЉE�}���  ~�   �I�E�E�}� ~:�U�H�E�H�@     H�4H��I��H�={������H��ЋE�Hc�H�E�H��  �E�H��0[A_]���UH��AWH����H�����I�vV      L؉}�H���������H�H�
�U�H�Ή�I��H�Ό������H���H��A_]���UH��AWSH�� ��H�����I�V      L�H�}�H�}� tj�E�    �?H���������H�H��E�Hc�H�E�H�� ��H�։�I��H�Ό������H��ЃE�H�E�H��I��H�"�������H��ЋU�9�w���H�� [A_]���UH��AWH���   ��L�����I�qU      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H���������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I�|T      M�H��8���H��0���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�H���������I�<M�׸    H�~�������L�������UH��AWH����H�����I��S      L�H�}�H�U�H��I��H�ة������H��ҐH��A_]���UH��AWH��(��H�����I��S      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H�W�������H��Ѹ    H��(A_]���UH��AWH��(��H�����I�-S      L�H�}�H�u�H�U�H�U�H�U�H�M�   H��I��H�W�������H����H�E�H�E�� < tH�E�H   H9E�sH�E�� <
u�H�E��  H�E�H;E�����H��(A_]���UH��AWSH��0��H�����I��R      L�H�}�H�uЉỦM�H�@	     H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H�W�������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H�@	     H�H�E�H�@	     �0H�@	     �D �}�u-�U�H�E�    H��I��H�&�������H���H�U�H��   �}�u+�U�H�E�    H��I��H�J�������H��Љ�H�EЉ�[�}�u,�U�H�E�    H��I��H�J�������H��Љ�H�E�f��)�U�H�E�    H��I��H�J�������H��Љ�H�EЈ�    H��0[A_]���UH��AWSH��0��H�����I��P      L�H�}�H�uЉỦM�H�@	     H�H�E�H�E�H   H�E�H�U�H�E�   H��I��H�W�������H����H�E�H�E�� < uH�E�� ��t
H�E�H;E�r�H�E�H;E�r/H�@	     H�H�E�H�@	     �0H�@	     �D �}�u'H�E�H��I��H���������H����Z�H�E�� �+�}�u%H�E�H��I��H���������H���fH~�H�U�H��    H��0[A_]���UH��SH��8��H�����I��O      L�H�}�H�u�H�U��E�    �E�    ��  �E�    �E�Hc�H�E�H�� ������%��  �E��E�Hc�H�E�H�� ������lu�E��E�   �E�Hc�H�E�H�� ����H���������H���	E�}��o  �E�H��    H��I  H�H�}I  H�>��H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H�`�������H�����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�H�E�H��H��H�Ŭ������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�g�������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�g�������H����  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��������H����?  H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�g�������H�����   H�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H�g�������H����jH�Eȋ ��/w$H�E�H�PH�Eȋ ��H�H�Uȋ�JH�Uȉ
�H�E�H�@H�HH�U�H�JH�0H�Eع
   �   H��H��������H������E��E�Hc�H�E�H�� ��������E�H��8[]���UH��H����H�����I�PK      L؉��E��E�    �E��S��%wa��H��    H�wF  H�H�lF  H�>���E�   �>�E�   �5�E�   �,�E�   �#�E�   ��E�   ��E�   ��E�������E�����UH��AWH���   ��L�����I��J      M�H�����H�����H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H�� ���H�����H�����H��H��M��H�H�������L��Љ�<�����<���H���   A_]���UH��AWH���   ��L�����I��I      M�H�����H��H���H��P���H��X���L��`���L��h�����t#)�p���)M�)U�)]�)e�)m�)u�)}�ǅ ���   ǅ$���0   H�EH��(���H��@���H��0���H���������I�H� H�� ���H�����H��H��M��H�H�������L��Љ�<�����<���H���   A_]���UH��H����H�����I��H      L؉}�H�u�H�}� u������w�}��u������jH�E��@#��tH�E��@#�P�H�E��P#H�E��@#H�U��J�    ��Љ�H�E�f�H�E�H�PH�E�� H��H�H�E�H�PH�E�H�@�U���E�����UH��AWSH����H�����I�H      L�H���������H�H� H��I��H�K!������H��ЉE�}��t+H���������H�H��E�H�։�I��H�/������H��ЋE�H��[A_]���UH��AWH��(��H�����I��G      L�H�}�H�u�H�U�H���������H�<I�ϸ    H�~�������H�������UH��H����H�����I�.G      L�H�}��	   H�E�H���r�����UH��SH����H�����I��F      L�H�}�H�}� u.H�@	     H�<H�Ƹ������H���H�@	     H��H�E�H��H�Ƹ������H���H�E�H��[]���UH��AWSH��0��H�����I�rF      L�H�}�H�u�H�E�H���������H�4H��I��H���������H���H�E�H�}� u
������   �E�    H�E�H��I��H�"�������H��ЉE܃}�`~	�E�   �$H�E�H�P+H�E�H��H��I��H�F~������H���H�E��@���H�E��PH�E�H��I��H�8�������H��ЋE�H��0[A_]���UH��H��0��H�����I�}E      L؉}�H�u�H�E�H�E��E܉E��E�    �}� y,H�E�H�PH�U�� -�}�   �u�E�����E���E��؉E�H�E�H�E�M�Hc�Hi�gfffH�� ��������)�����)��ʉЍH0H�E�H�PH�U�ʈ�E�Hc�Hi�gfffH�� ����)ЉE�}� u��}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWSH��@��H�����I�3D      L�H�}�H�u��U�H�}� u#H�E�H�E�H�E�H�PH�U�� 0H�E��  �  H�E�H�E؋E�Hc�H�E�H�H�E��3H�E؃��E�H�m��}�	~�7   ��0   �U��H�m���H�E�H�E�H;E�wËE�Hc�H�E�H��  H�E�H�E��E�    �8H�E�� <0uH�E��"H�U�H�E�H��H��I��H�F~������H�����E��E�;E�|�H�E�H�E�H�E�H��I��H�"�������H��Љ�H�E؋E�H�U�)Љ�H�M�H�E�HȾ    H��I��H��{������H���H��@[A_]���UH��AWH����H�����I��B      L؉}�U�    ��I��H��O������H���H��A_]���UH��AWH����H�����I�rB      L؉}�u�U��U��I��H�3�������H���H��A_]���UH��AWH����H�����I�#B      L�H�}�H�U�H��I��H��R������H��ҐH��A_]���UH��AWH����H�����I��A      L�H�}�u�M�H�U��H��I��H��T������H���H��A_]���UH��H����H�����I��A      L؉}�u�E��}�E��E��}�ЉE��}� x�E���y�E����E��E�+E�E��!�}� y�E���~�E����E��U��E�ЉE�H�E�����UH��H�� ��H�����I��@      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H�� ��H�����I�T@      L�H�}�H�u�H�E�H�H�}�H�E�H�E�H�H�}�H��H�E�H�}� x#H�E�H��yH�E�H��H�E�H�E�H+E�H�E��+H�}� y$H�E�H��~H�E�H��H�E�H�U�H�E�H�H�E�H�E�H�U�����UH��H��H��H�����I��?      L�H�}�H�u��U�H�E�H�E�H�E�H�PH�U�� ���E�E���H���������H�H������ ��uǃ}�-u�E�   H�E�H�PH�U�� ���E��"�E�    �}�+uH�E�H�PH�U�� ���E�}� t�}�u9�}�0u3H�E�� <xtH�E�� <XuH�E�H��� ���E�H�E��E�   �}� u�}�0u�   ��
   �E��}� t	H��   ������H�E�E�Hc�H�E�H�H��H�ЉE؋E�Hc�H�E�H�H��H�E�}� t�}� ~�E�)E�H�E��]�H�E�    �E�    �E���H���������H�H��������t�m�0�[�E���H���������H�H���������5  �E���H���������H�H��������t�7   ��W   )E�E�;E���   �}� ��   �}� tgH�E�H;E�|H�E�H;E�u0�E�;E�~(�E�����H�E�   �H���������H�� �����   �E�   �E�H�H�U�H��H�E��E�H�H)E��eH�E�H;E�H�E�H;E�u-�E�;E�~%�E�����H�E����H���������H�� �����$�E�   �E�H�H�U�H��H�E��E�H�HE���H�E�H�PH�U�� ���E��y������H�}� t�}� t
H�E�H���H�E�H�U�H�H�E�����UH��AWH����H�����I�v<      L�H�}�H�M�
   �    H��I��H�J�������H���H��A_]���UH��AWH����H�����I�!<      L�H�}�H�M�
   �    H��I��H�J�������H���H��A_]���UH��AWAVAUATSH����H�����I��;      L�H�}�H�uȉU�L�eп    L��L�`� �؉���H���������H�H������ ��uЃ�-u�   L��L�`� �����+uL��L�`� �؃}� t�}�u-��0u(A�$<xt	A�$<XuI�D$� ��I���E�   �}� u��0u�   ��
   �EċE�Hc������    H��I�ǋE�Hc������    H��H�Љ�A�    A�    ����H���������H�H��������t��0�T����H���������H�H��������tz����H���������H�H��������t�7   ��W   )�;]�}GE��x
M9�wM9�u��9�~A������A�   �E�H�L��Hc�I�L��L�`� ���;������E��yA�����H���������H�� "   �	����tI��H�}� tE��tI�D$��H�E�H�U�H�L��H��[A\A]A^A_]���UH��H����H�����I��9      L؉}��   �   ���r����UH��AWSH����H�����I�H9      L�H�}�H�E�H���������H�4H��I��H��}������H��Ѕ�uH���������H�H� ��    H��[A_]���UH��AUATSH�� ��H�����I��8      L�H�}�H�u�H��	     ��E�L�e�H�]�E�,$L��L�`��H��H�XD�(�m��}� uې�H�� [A\A]]���UH��H��8��H�����I�Y8      L�H�}�H�u�H�U�H��	     ��E�H�E�H�E�H�E�H�E�H�E�H�E�H�E�� ���E�H�E�H�PH�U�H�U���H�E�H�PH�U�H�U���H�E�H�PH�U��U���m��}� u�������UH��SH��H��H�����I��7      L�H�}�H�u�H��	     ��E�H�E�H+E��EȋE�9E���  �E�����EȺ    ��E��EȋU�H�E�H�H�E�H�E�H�E�H�E�H�E�E�H�H��H��H�E�H�H�E�H�E�H;E�sjH��	     H�H�U�H�E�H��H���щEă}� u/�E�H�H��HE�H�U�H�E�H��H��H� �������H�����  �}� y�E�H�HE���  �H�E�H;E���   H��	     H�H�U�H�E�H��H���щEă}� u)�E�H�HE�H�U�H�E�H��H��H� �������H���뢃}� ��   H�E�H;E�uA�E�H�HE�H�U�H�M�H�E�H��H��H���������H��ЋE�H�HE�H�E�H�E��M���H�U�H�E�H��H��H� �������H��ЋE�H�H��HE��E�H�HE���   �E�H�H��HE�����H�E�H;E���   H�E�H+E�H��H�E�H+E�H9�|4�E�Hc�H�E�H�H�E�H��H��H�I�������H���H�E�H�E������H�U�H�E�H��H��H�I�������H��ЋE�Hc�H�E�H�H�E������E�H�H��HE�H�U�H�M�H�E�H��H��H���������H��ЋE�H�H��HE�H�E�H�E������H��H[]���UH��H�� ��H�����I��4      L�H�}��u�U�H�M�H��	     H�U�H��U�H��	     ��U��U���H�U�H�H�U�H��H��H�I�������H��А����UH��AWH����H�����I�64      L�H�}�H���������H�<I�׸    H�~�������H��Ѹ����H��A_]���UH��H��@��H�����I��3      L�H�}�H�u�H�U�H�U��H�E�H�U����H���������H�Hc���҃� ��u��E�    H�U���҃�+t��-u�E�   H�E�H�����������E��E�    �E�    �E�    �;�M�H�����������Y�H�U���҃�0�*��X��E�H�E��E�H�U����H���������H�Hc���҃���u�H�U����.uuH�E��?�M�H�����������Y�H�U���҃�0�*��X��E�H�E��E��E�H�U����H���������H�Hc���҃���u��U�)U�}� uH���������f���  �}� t�E�H���������f(fW��E�H�U����etH�U����E��   �E�    H�E�H�U���҃�+t��-u�E�   H�E��E�    �%�M܉����҉�H�U���҃�0ʉU�H�E�H�U����H���������H�Hc���҃���u��}� t�U�)U���U�U�}����|	�}�   ~H� ���������   H�����������E��E�E܃}� yF�]��A�E܃���t&�}� y�E��^E��E���E��YE��E��}��E��Y��E��}� u�H�}� tH�E�H�U�H��E�����UH��H����H�����I��0      L؉}�H�E�   �E�    �H�U�H��H��H�H�H�E��E��E�;E�|�H�E�����UH��AWSH��@��H�����I�E0      L��E�H�}��u�H�}� u	H�E��  H�E�H�E�H���������f��f/E�v,H�E�H�PH�U�� -�E�H� �������f(fW��E��E�H��������f/s�E��H,�H�E��/�E�H����������\��H,�H�E�H�       �H1E�H�E�H�E�H�E�H��x�H*��H��H���H	��H*��X��M��\�f(��EȋE���H�M�������H���H��x�H*��H��H���H	��H*��X��YE�H��������f/s�H,�H�E��*H����������\��H,�H�E�H�       �H1E�H�E�H�E�H�M�H�U�H�E�H���������H�43H��I�߸    I���������I�A��H�E�H��@[A_]���UH��AWH����H�����I�[.      L�H�}�H�U�    H��I��H��������H���H��A_]���UH��AWH����H�����I�.      L�H�}�H�u�H�M�H�U�H��H��I��H��������H����Z�H��A_]���UH��AWH��(��H�����I��-      L�H�}�H�u�H�M�H�U�H��H��I��H��������H����E��E�H��(A_]���UH��H����H�����I�U-      L؉}��E����3E�)�����UH��H��@��H�����I�!-      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�    H�}� y>H�E�H�PH�U�� -H�       �H9E�uH��������H�E�H�E��H�E�H��H�E�H�E�H�E�H�M�H�gfffffffH��H��H��H��H��?H)�H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U��ʈH�M�H�gfffffffH��H��H��H��H��?H)�H��H�E�H�}� u�H�}� tH�E�� ����H�E��H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U߈H�E�H;E�w�H�E�����UH��AWH��8��H�����I��+      L�H�}�H�uЉU�H�U�H�U�H�}� yH�U�H�JH�M��-H�]�H�U�H�U��}�u$H�M�H�u�   H��I��H���������H����H�M�H�U�H��H��H���������H���H�E�H��8A_]���UH��H��0��H�����I��*      L�H�}�H�u�H�E�H�E�H�E�H�E�H�E�H�E�H�M�H���������H��H��H��H��H��H�H�H)�H�ʉЍH0H�E�H�PH�U�ʈH�E�H���������H��H��H��H�E�H�}� u�H�E�H�P�H�U��  �1H�E�� �E�H�E�H�PH�U�H�U���H�E�H�P�H�U��U�H�E�H;E�w�H�E�����UH��AWH��8��H�����I�*      L�H�}�H�uЉU�H�U�H�U�H�U�H�U��}�u$H�u�H�M�   H��I��H���������H����H�M�H�U�H��H��H���������H���H�E�H��8A_]���UH��H����H�����I�n)      L؉}������UH����H�����I�H)      Lظ   ]���UH��H����H�����I�)      L�H�}��    ����UH��H����H�����I��(      L�H�}�H���������H�H� ����UH��H����H�����I��(      L�H�}�H���������H�H� ����UH��H�� ��H�����I�x(      L�H�}��u�H�U�H�M�    ����UH����H�����I�B(      Lظ    ]���UH��H����H�����I�(      L��E�H��������f������UH��H����H�����I��'      L��E�H��������f������UH��H����H�����I��'      L��E��}�H��������f������UH��H����H�����I�i'      L��E�H�}�H��������f������UH��H����H�����I�,'      L��E��M�H��������f������UH��H��(��H�����I��&      L��E��M��E��U��U��E��E��E������������������������������]��E�����UH��H����H�����I��&      L��E����E����]��E�����UH��H����H�����I�E&      L��E�H� �������f������UH��H����H�����I�&      L��E�H�(�������f������UH��H����H�����I��%      L��E�H�0�������f������UH��H����H�����I��%      L��E�H�8���������E��E�����UH��H����H�����I�V%      L��E�H�@�������f������UH��H����H�����I�%      L��E�H�H�������f������UH��H����H�����I��$      L��E�H�P�������f������UH��H����H�����I��$      L��E�H�X�������f������UH��AWH����H�����I�p$      L��E��E�H�`�������H�f(�fHn�I��H��������H���H��A_]���UH��H����H�����I�$      L؉}�H�u�    ����UH��AWH����H�����I��#      Lډ}�H�u�H�h�������H�<I�׸    H�~�������H�������UH��AWH��(��H�����I��#      Lى}�H�u�H�U�H�y�������H�<I�ϸ    H�~�������H�������UH��AWSH�� ��H�����I�0#      L�H�}�H���������H�<I�߸    H�~�������H����E�    �.�E�H�H��    H�E�HЋ ��I��H�|�������H��ЃE��}�?~̸����H�� [A_]���UH��AWH����H�����I��"      L�H�}�u�H���������H�<I�׸    H�~�������H�����f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     f.�     fD                                                                      ~ � � � � � � � � ~             ~ � � � � � � � � ~                 l � � � � | 8                   8 | � | 8                   < < � � �   <                < ~ � � ~   <                      < <              � � � � � � � � � � � � � � � �           < f B B f <           � � � � � � � � � � � � � � � �        2 x � � � � x             < f f f f <  ~               ? 3 ? 0 0 0 0 p � �              c  c c c c g � � �               � < � < �             � � � � � � � � � � �               > � >                  < ~    ~ <                f f f f f f f   f f              � � � {                | � ` 8 l � � l 8  � |                       � � � �              < ~    ~ <  ~              < ~                           ~ <                      �                         0 ` � ` 0                         � � � �                       ( l � l (                      8 8 | | � �                   � � | | 8 8                                                 < < <                  f f f $                             l l � l l l � l l           | � � � |   � � |               � �   0 ` � �             8 l l 8 v � � � � v           0 0 0 `                             0 0 0 0 0 0               0         0                   f < � < f                         ~                                    0                     �                                                           0 ` � �             8 l � � � � � � l 8              8 x       ~             | �    0 ` � � �             | �   <    � |               < l � �                 � � � � �    � |             8 ` � � � � � � � |             � �     0 0 0 0             | � � � | � � � � |             | � � � ~     x                                                       0                  0 ` 0                      ~     ~                     ` 0      0 `             | � �                       | � � � � � � � |              8 l � � � � � � �             � f f f | f f f f �             < f � � � � � � f <             � l f f f f f f l �             � f b h x h ` b f �             � f b h x h ` ` ` �             < f � � � � � � f :             � � � � � � � � � �             <         <                   � � � x             � f f l x x l f f �             � ` ` ` ` ` ` b f �             � � � � � � � � � �             � � � � � � � � � �             | � � � � � � � � |             � f f f | ` ` ` ` �             | � � � � � � � � |           � f f f | l f f f �             | � � ` 8   � � |             ~ ~ Z       <             � � � � � � � � � |             � � � � � � � l 8              � � � � � � � � � l             � � l | 8 8 | l � �             f f f f <     <             � � �   0 ` � � �             < 0 0 0 0 0 0 0 0 <               � � � p 8                 <         <          8 l �                                                   �       0                                     x  | � � � v             � ` ` x l f f f f |                   | � � � � � |                < l � � � � v                   | � � � � � |              6 2 0 x 0 0 0 0 x                   v � � � � � |  � x       � ` ` l v f f f f �                 8      <                        f f <       � ` ` f l x x l f �             8         <                   � � � � � � �                   � f f f f f f                   | � � � � � |                   � f f f f f | ` ` �             v � � � � � |                � v f ` ` ` �                   | � ` 8  � |              0 0 � 0 0 0 0 6                    � � � � � � v                   � � � � � l 8                   � � � � � � l                   � l 8 8 8 l �                   � � � � � � ~   �             � �  0 ` � �                 p                                        p         p                       v �                        8 l � � � �                               ��� ��� ~~~                                 uuu ��� ��� ���                                 ��� ��� ��� ��� ;;;                          ��� ��� ~~~ ��� ���                         ��� ��� ���     ��� ���                         ��� ���      ��� ��� ppp                 @@@ ��� ���         III ��� ���                 ��� ��� ��� ��� ��� ��� ��� ���                 ��� ���                 zzz ��� ���         ``` ��� ���                     ��� ���         ��� ��� MMM                     ��� ��� bbb     ��� ���                         ||| ��� ���      ��C                        Usage: %s <input.jpg> [<output.ppm>]
 rb        Error opening the input file.
  Error decoding the input file.
 nanojpeg_out.ppm nanojpeg_out.pgm w+b   Error opening the output file.
 P%d
%d %d
255
                           	
 !(0)"#*1892+$%,3:;4-&'.5<=6/7>?�#������l$������l$������l$������$������l$������l$������l$������l$������l$������l$������l$������l$������l$������l$������l$������l$������l$������l$������l$������l$������l$������l$������l$������l$������l$������H$������$$������l$������6$������Entrada maior que o limite
 Erro ao criar o arquivo "%s"
       Error ao criar o arquivo "%s", atingio o limite de arquivos na entrada de directorio
   Panic: __malloc, sem espaco na tabela de alocacao
      panic: realoc sem espaco, %lx size = %d %d
 PWD BitMAP error
 Not suport BitMAP 4-bit Not suport BitMAP > 8-bit strerrorr
      (((((�AAAAAABBBBBB                                �Dubug: %s %x %x
        (null)  ڣ���������������������E����������������������L�������L�������ڣ������ڣ������ڣ������ڣ������ڣ������ڣ������ڣ������ڣ������ڣ������ڣ������ڣ���������������������l���������������������<�������r�������r�������r�������r�������W�������r�������r�������r�������r�������r�������r�������r�������r�������r�������r�������3�������E�������r�������i�������`�������r�������E�������r�������r�������r�������r�������r�������r�������r�������r�������r�������<�������r�������N�������r�������r�������W�������(null) %        ~���������������6����������������������G�����������������������~�������~�������~�������~�������~�������~�������~�������~�������~�������~�������~���������������a��������������ë������ë�������������H�������H�������H�������H�������-�������H�������H�������H�������H�������H�������H�������H�������H�������H�������H�������	��������������H�������?�������6�������H��������������H�������H�������H�������H�������H�������H�������H�������H�������H��������������H�������$�������H�������H�������-�������panic: sscanf()
        չ���������������������S���������������չ������+�������+�������չ������չ������չ������չ������չ������չ������չ������չ������չ������չ������չ���������������������չ������l�������l���������������ٹ������ٹ������ٹ������ٹ��������������ٹ������ٹ������ٹ������ٹ������ٹ������ٹ������ٹ������ٹ������ٹ������ٹ����������������������ٹ������й������ǹ������ٹ��������������ٹ������ٹ������ٹ������ٹ������ٹ������ٹ������ٹ������ٹ������ٹ��������������ٹ��������������ٹ������ٹ��������������panic: freopen()
 r+ PWD call system funtion error. 
                 $@       �        %lu.%lu                �              �C                                                                        �_�
�@panic: signal()
 panic: sigaction()
 panic: setjmp()  panic: longjmp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    F
 �     �     �   �N
 �   F
 �   �N
 �      �   8F
 �      �   �5 �   HF
 �   hF
 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          zR x�  ,      @����   E�CG����B�A�       0   L   �����   E�CK����u�B�B�B�A�      �   H���I    E�C@�    �   q����   E�C��$   �   ����   E�CE���A�      �   �����   E�C��      9����    E�CE�q�A�    ,  ����_    E�CE�P�A�   P  ����M    E�CD�    p  �����    E�C��    �  ����I    E�C@�     �  �����    E�CA���A�    �  Y���U    E�CA�J�A�(   �  ����	   E�CG����B�A�   (   $  g����   E�CG����B�A�   $   P  ����c   E�CE�T�A�       x  ����    E�CA���A�$   �  ����"   E�CE��A�   (   �  �����   E�CG����B�A�   $   �  L����   E�CE���A�   ,     �����   E�CI�����B�B�A�   (   H  +����   E�CG����B�A�   4   t  ����p   E�CM�����Q�B�B�B�B�A�       �  ��Y    E�CF�I�A�$   �  =��    E�CG����B�A�$   �  ���   E�CE���A�         ���0    E�Cg�     @  ���0    E�Cg�     `  ���9    E�Cp�     �  ���X    E�CO�     �  ��R    E�CI�     (   �  5��Z   E�CG��G�B�A�      �  c��   E�C�     a���    E�C��    0  ����    E�C��     P  r��p    E�CF�`�A�$   t  ����    E�CG����B�A�$   �  }	��r    E�CG��_�B�A�(   �  �	��   E�CG��	�B�A�   $   �  ����   E�CF���A�         ^���    E�CE���A�    <  ����    E�CE���A�   `  ����    E�C��    �  I��A    E�Cx�      �  j��i    E�C`�        �  ���U    E�CL�    �  ���U    E�CL�      ��i    E�C`�    $  b��g    E�C^�    D  ����    E�C�� $   d  p���   E�CE�{�A�      �  ���9    E�Cp�  $   �  ����    E�CG����B�A�   �  ���^    E�CU� (   �  ���   E�CG���B�A�   (      ����   E�CG����B�A�   (   L  q��]   E�CG��J�B�A�   (   x  ���   E�CG��l�B�A�   (   �  ���D   E�CJ��.�B�A�   (   �  $��:   E�CG��'�B�A�   $   �  %��    E�CG����B�A�   $	  �%���    E�C��    D	  �&���    E�C�� (   d	  ['���   E�CJ����B�A�   (   �	  +��i   E�CG��V�B�A�   (   �	  [.��H   E�CG��5�B�A�   (   �	  w0��e   E�CJ��O�B�A�      
  �4��a    E�CX�    4
  �4��9    E�Cp�      T
  
5���    E�CF�w�A�(   x
  m5��'   E�CG���B�A�   $   �
  h8��   E�CE���A�   $   �
  A:���   E�CF���A�      �
  �;��    E�C��      �<���    E�C�� (   4  _=��O   E�CG��<�B�A�   $   `  �>���    E�CG����B�A�(   �  F?��C   E�CG��0�B�A�      �  ]A��k    E�Cb� $   �  �A���    E�CG����B�A�   �  hB���    E�C�� $     �B��   E�CE��A�   $   D  �C���    E�CG����B�A�$   l  RD���    E�CG����B�A�(   �  �D���   E�CG����B�A�   (   �  oF��j   E�CG��W�B�A�       �  �G���    E�CE���� (     EH��   E�CG���B�A�       <  8I���    E�CE���� (   `  �I���   E�CG��q�B�A�   $   �  (N��   E�CG����B�A�   �  O��9    E�Cp�     �   O��+    E�Cb�     �  +O���    E�C��       �O���   E�CE����   8  :R��I    E�C@�     X  cR��u    E�CE�f�A�(   |  �R���   E�CG����B�A�   (   �  jU���   E�CG����B�A�   $   �  !X���    E�CG����B�A�,   �  �X��2   E�CG���B�A�          ,  �[���    E�C��    L  M\��w    E�Cn�    l  �\��b    E�CY� $   �  �\���    E�CG����B�A�$   �  y]��z    E�CG��g�B�A�   �  �]��a    E�CX�    �  ^���    E�C��      �^��{    E�Cr� $   <  �^��+   E�CF��A�      d  �_��6   E�C-�   �  �`��L    E�CC� $   �  &a���    E�CG����B�A�   �  �a���    E�Cw�    �  &b��}    E�Ct� $     �b��r    E�CF�b�A�    $   4  �b���    E�CF���A�       \  8c���    E�C��    |  �c��3   E�C*�   �  �d��7   E�C.�   �  �e��W    E�CN� $   �  6f���    E�CG����B�A�$     �f���    E�CG����B�A�   ,  g���    E�C�� $   L  �g��V    E�CF�F�A�       t  �g��P    E�CF�       �  h��U    E�CL�    �  Sh��U    E�CL� $   �  �h���    E�CG����B�A�$   �  i���    E�CG����B�A�$   $  pi��K    E�CF�{�A�     $   L  �i��K    E�CF�{�A�     $   t  �i��S    E�CF�C�A�    $   �  �i���    E�CG����B�A�$   �  Qj��S    E�CF�C�A�    $   �  |j��K    E�CF�{�A�     ,     �j��[   E�CG��H�B�A�       $   D  �k���    E�CG����B�A�$   l  Fl��]    E�CF�M�A�    $   �  {l��]    E�CF�M�A�    $   �  �l��K    E�CF�{�A�     $   �  �l��L    E�CF�|�A�     $     �l��Y    E�CF�I�A�       4  (m��Y    E�CP� $   T  am��K    E�CF�{�A�     (   |  �m���   E�CJ��{�B�A�       �  �u���    E�C��     $   �  ov���    E�CI���A�       �  2w��l    E�Cc� (     ~w���   E�CJ����B�A�       @  '����    E�C��     $   d  ����   E�CI���A�    $   �  �����    E�CI���A�    $   �  K����    E�CG����B�A�$   �  ����\    E�CF�L�A�    $     0����    E�CG����B�A�$   ,  �����    E�CI���A�       T  {����    E�CI�    $   t  ����L    E�CF�|�A�         �   ���e    E�CF�U�A�    �  a����    E�CF���A�(   �  ߅���   E�CG����B�A�   (     W���=   E�CG��*�B�A�   $   <  h���\   E�CE�M�A�      d  �����    E�C�� $   �  &����    E�CI���A�    $   �  ����    E�CI���A�       �  �����    E�C�� $   �  H����    E�CG��z�B�A�     ����Y    E�CF�       <  ���9    E�Cp�  $   \  �����    E�CE�q�A�    $   �  W����    E�CG����B�A�   �  '���G   E�C>�,   �  N���u   E�CG��b�B�A�       $   �  ����M    E�CF�}�A�     $   $  ����O    E�CF��A�     $   L  ߓ��L    E�CF�|�A�     $   t  ���S    E�CF�C�A�       �  .����    E�C�    �  �����    E�C��    �   ����    E�C��    �  ����2   E�C)�$     ����U    E�CF�E�A�    $   D  ���U    E�CF�E�A�    4   l  ���L   E�CM�����-�B�B�B�B�A�      �  *���7    E�C       $   �  A���w    E�CG��d�B�A�(   �  ����{    E�CI���d�B�B�A�     ߛ���    E�C�� $   8  m����   E�CE���A�       `  7����    E�Cx�     $   �  ����\    E�CF�L�A�       �  ȟ��5   E�C,�   �  ݢ��_    E�CV� ,   �  ����   E�CG����B�A�       $     פ��P    E�CF�@�A�    $   D  ����Z    E�CF�J�A�    $   l  1���^    E�CF�N�A�       �  g���4    E�Ck�     �  {���v   E�Cm�$   �  Ѧ���    E�CF���A�       �  X����    E�C�� $     1����    E�CF���A�       D  ����*    E�Ca�     d  ����'    E�C^�     �  ����/    E�Cf�     �  ����;    E�Cr�     �  ٨��;    E�Cr�     �  ����:    E�Cq�       ���'    E�C^�     $  ���9    E�Cp�     D  .���9    E�Cp�     d  G���<    E�Cs�     �  c���=    E�Ct�     �  ����>    E�Cu�     �  ����n    E�Ce�    �  ���;    E�Cr�        ���9    E�Cp�     $    ���9    E�Cp�     D   9���9    E�Cp�     d   R���D    E�C{�     �   v���9    E�Cp�     �   ����9    E�Cp�     �   ����9    E�Cp�     �   ����9    E�Cp�  $   !  ڪ��a    E�CF�Q�A�       ,!  ���2    E�Ci�     L!  %���T    E�CF�   h!  ]���X    E�CF�$   �!  �����    E�CG����B�A�   �!  ���T    E�CF�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            GCC: (Ubuntu 9.3.0-17ubuntu1~20.04) 9.3.0                                        �                    �                  @ �                 `@ �                 �@ �                  P
 �                                     ��                     ��_ cole _             ��                )        �                    �           0    ��                7    ��                B     �@ �   �     E     `3 �   @       J     �,  �   �      U     q0  �   �       \     l1  �   �       k     pC	 �          w     D>  �   "      �      �2 �           �      �2 �           �      �2 �           �      �2 �           �      �2 �           �      3 �           �      3 �           �      3 �           �      83 �           �    ��                �    ��                �      �4 �           �      �4 �           �      �4 �           [   ��                �     �C	 �          �      (5 �           �      `5 �           �    ��                �    ��                �      �5 �           �    ��                �    ��                �    ��                �    ��                �      �5 �           �      �5 �           �      �5 �           �    ��                �    ��                   ��                   ��                   ��                #   ��                0   ��                9   ��                B   ��                K   ��                T   ��                ^   ��                g   ��                p   ��                ~   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �    �C	 �          �   ��                �   ��                �   ��                �   ��                �   ��                �      �5 �           �   ��                   ��                   ��                   ��                �      �6 �               ��                (   ��                1   ��                ;   ��                C   ��                :   ��                B   ��                J   ��                R   ��                Z   ��                b   ��                k   ��                t   ��                }   ��                �   ��                �   ��                �   ��                �    ��  �   �       �      �6 �           �   ��                �   ��                �    k�  �   �       �      �8 �           �      �8 �           �   ��                �   ��                �   ��                �    �C	 �          �   ��                S   ��                �   ��                �   ��                �      �: �           �   ��                �   ��                �    ��  �   e       &    %�  �   �       �    ��  �   �      �    �C
 �          �    k�  �   =          �D
 �          �    �  �   �       �   ��                �   ��                   ��                   ��                   ��                �      �< �           (   ��                1    �E
 �   `       9   ��                �      
= �           B   ��                I   ��                Q   ��                Z   ��                c   ��                j   ��                v   ��                u   ��                t   ��                |   ��                �   ��                �   ��                �   ��                �   ��                �   ��                �      = �           �   ��                �     F
 �          �    F
 �          �    � �   {       �    � �   �       �    � �   �      �   ��                �      = �           �   ��                �      0= �           �      8= �           �      @= �           �   ��                �    � �   _       �      X= �           �      `= �           �      p= �           �      P= �           �   ��                �   ��                   ��                   ��                   ��                   ��                #   ��                $   ��                +   ��                L   ��                3   ��                <   ��                H   ��                S   ��                [   ��                �      x= �           b   ��                h   ��                o   ��                �      �= �           v   ��                �      �= �           }   ��                �      �= �           ~   ��                �      �= �           p   ��                �      �= �           w   ��                �      �= �           �   ��                �      �= �           �   ��                �      �= �           �   ��                �      �= �           �   ��                �   ��                �      �= �           �      �= �           �   ��                �      �= �           �      �= �                ��                �    `@ �           �    � �   T       �    �k  �         �    ��  �   \       �    1<  �   c      �    ��  �   �       �    ��  �   {           v �   9           � �   ;           ! �   �           ��  �   �           �j  �   �       '    ��  �   7      0    �T  �   Y       C    ��  �   �       7    F
 �          >    ��  �   �      G    ��  �   �       N      �           V    V  �   �      _    �/  �   _       �    �  �   �       i      �           n    f�  �   P       w    X �   �       ~    �N
 �          �    N�  �   �       �    �  �   �       �    F
 �          �    �  �   �      �    1 �   U       �    ��  �   u       �    	 �   w       �    � �   9       �    �X  �   0       �    �N
 �          �    p �   9       �    � �   ^       �    `2 �          �    � �   �       0    ��  �   �       �    ��  �   [      �    �|  �   :      �      �   �           �2  �   	      v
    ��  �   �           ��  �   w       !    #1  �   I       ,    #�  �   �       ;    12  �   U       H    �  �   �      P    t�  �   L       W    3 �   v      �    8�  �   �       ^    ��  �   U       f     �   \       m    `�  �   Y       r    ��  �   M       y    p�  �   K       !
     F
 �          �    �F
 �          �    ��  �   �      �    � �   <       �    �  �   �       �    � �   L      �    ��  �   G      �    (F
 �          �    W[  �         �    �o  �   ]      �       �   �       �    ��  �   K       �       �           �    ��  �   �          4�  �   �           P
 �               �Y  �   Z          �  �   �       $    �e  �   A       +    ��  �   �       7    @B  �   �      D    շ  �   2      K    ;d  �   �       S    �  �   2      Z    0F
 �          _    ��  �   �       f    6^  �   �       n    �  �   �       v    Q �   �       {    ��  �   O       �    x �   5      �    f  �   i       �    � �   P       �    wK  �   �      B    ?�  �   �       �    �d  �   �       �    1�  �   z       �    �m  �   �           �
 �           �    `�  �   �       �    �  �   Y       �    �%  �   I       �    )�  �   9       �    À  �   �      �     �   �      -    7 �   9       �    8F
 �          �       �          k
    �@ �               �N
 �                 �               @F
 �               �
 �           #    �  �   �       *    bj  �   9       4    �g  �   g       �
    � �   D       �	     �   '       B    ( �   >       H    u �   T       O    �  �   V       W    ��  �   �       _    �f  �   U       l    E/  �   �       w    ��  �         �    �X  �   0       �    f �   n       �    �  �   }       �    h�  �   �       �    v�  �   �       �    = �   9       �    �F
 �          �    {�  �   S       �    3�  �   j      �    �(  �   �      �    �  �   k       �    r  �         l
    �@ �           �    &  �   �      	    ��  �   W       	    �  �   H      	    �  �   �       	    ��  �   �       !	    ��  �   �       -	    ~  �          8	    ��  �          C	    � �   X       M	    zc  �   �       T	    �  �   �       e	    ��  �   ]       k	    �5 �          r	    �u  �   D      |	    �N
 �          �	    �h  �   �      �	    ��  �   �       �	    $0  �   M       �	    Y  �   9       �	    �  �   �       
       �           �	    &�  �   9       �	    � �   ;       �	    �  �   b       �	    HF
 �          �	    <"  �   �      �	    �=  �   �       �	    ��  �   K       �	    � �   *       �	    ��  �   K       �	    �9  �   �      
    @�  �   �           7 �   /       
    _  �   r       
       �           
    PF
 �          2    _�  �   �       �    � �   a       (
    �  �         �
    .�  �   S       1
    ��  �   +       �    �a  �   �      ?
    ]  �   �       G
    *�  �   l           �_  �         Q
    �  �   �       q
    � �   9       X
    v�  �   I       ^
    c�  �   e      j
    �@ �           p
     �   9       u
    l�  �   K       ?    �  �         {
    Y�  �         �
    G �   Z       �
    L�  �   6      �
    � �   9       �
    � �   �       �
    C �   2       1    ��  �   �       �
    XF
 �          �
    ��  �   i      �
    ��  �   �       �
    u\  �   �       �
    �  �   '          V�  �   �       
       �           �
    `F
 �          �
    �  �   S       �
    �]  �   p       �
     0 �   @      �
    N   �           �
    Қ  �   C      
    � �   :           �  �   u             �   �           �  �   ]       &    hF
 �               �
 �           /    ��  �   \      7    ��  �   L       >    ��  �   Y       F    f?  �   �      �       �           T    ��  �   �       ^    � �   7       c    �F  �   �      o    pF
 �          v    �Y  �   R       �    Ȏ  �   a       �    � �   U       �    SY  �   X       �    ��  �         �    b�  �   �       (    4�  �   �      �    !g  �   i       �    f �   ;       �    U�  �   3      �    `   �   �      �    x�  �   �       �    ��  �   L       �       �           �    �  �   U       �    ��  �   9       �    U  �          �    �g  �   �            �   '       �       �           
    �k  �   ^           ��  �   �           � �   4           ��  �   a       &    �  �   �       ,    H �   9       1    !�  �   +      ;    � �   =       A    �  �   �      J    ��  �   r       R    wf  �   U       ^    /�  �   L       c    ��  �   O      k    HP  �   p       lib/setup.asm HEADER_MAGIC HEADER_FLAGS header crt0.c nanojpeg.c nj njZZ njShowBits njSkip njDecodeLength counts.1861 njGetVLC .LC0 .LC1 .LC2 .LC3 .LC4 .LC5 .LC6 .LC7 .LC8 file.c cfs.c alloc_spin_lock pipe.c path.c gui.c font8x16.c window.c bmp.c font.c border.c memcmp.c memcpy.c memset.c strcasecmp.c strcat.c strchr.c strcmp.c strcpy.c strcspn.c string.c strlen.c strncasecmp.c strncmp.c strncpy.c strpbrk.c strrchr.c strsep.c strspn.c strtok.c last.1481 strstr.c strdup.c memmove.c strcoll.c strerror.c ctype.c tolower.c toupper.c stdio.c fopen.c fclose.c fflush.c fputc.c fgetc.c fgets.c fputs.c fread.c fwrite.c remove.c rewind.c fseek.c feof.c ftell.c vfprintf.c vf vsprintf.c vsnprintf.c sn_buf putchar.c sscanf.c perror.c vfscanf.c character _buf.1638 fvalue _buf.1650 ungetc.c getchar.c freopen.c tmpnam.c _tmpnam rename.c itoa.c i2hex.c malloc.c calloc.c free.c realloc.c lldiv.c strtol.c atoi.c atol.c strtoul.c exit.c getenv.c qsort.c qscmp qses qsexc qstexc qs1 system.c strtod.c ftoa.c _precision atof.c strtof.c strtold.c abs.c ltoa.c utoa.c srand.c errno.c gmtime.c localtime.c strftime.c clock.c math.c pow.c sqrt.c atan.c acos.c asin.c floor.c ceil.c exp.c locale.c signal.c setjmp.c _GLOBAL_OFFSET_TABLE_ longjmp read_directory_blk njDecodeDQT drawstring strcpy log sqrt setjmp put clean_blk_enter strtok_r njInit stdout vsprintf ungetc pwd_ptr njDecode njGetBits argv strerror utoa_r __m_i memmove __tm __realloc_r atol __window_puts getenv ceil njGetHeight errno floor strtold _infinity qsort fgets file_update file_read_block njDecodeSOF memcpy njDecode16 __window_clear njSkipMarker BitMAP2 perror ltoa_r tolower system feof malloc remove fs_directory __window_putchar ldexp vsnprintf strtoul itoa __pipe__ stdgetc_r update_directory_entry _drawline fflush argc drawrect BitMAP eh_frame stdputc_r upath tell_r strncasecmp njDecodeScan border write_r strtol user rename flush_r strrchr utoa calloc strtod rewind_r atof njUpsampleV seek_r strcat read_directory_entry debug_o fseek njClip __free_block_r open_dir ftoa stdin font8x16 __m_c _start obj_list __end strstr write_blk get_file_name atan2 signal strcoll strncmp write_sector njSkipBits draw_char_transparent njGetWidth pow strncpy put_pixel strcasecmp log10 _BLK_ realloc drawchar njColIDCT path_count open_file_r njRowIDCT strtok remove_blk memcmp sscanf getfilename file_close pipe_write sigaction read_r file_write_block fread _ctype open_file addr search_blk_null strdup njByteAlign njIsColor fopen sysgettmpnam localtime memset pwd main njDecodeDRI ftell srand fclose njDecodeDHT getchar close_r __data ptr_mouse2 __free_r update_window getkeyw _vsputs_r strcmp color remove_file __bss atan fgetc drawchar_trans strtof strcspn asin ltoa setlocale stderr create_file strsep getkey __malloc_r mouse fputc open_r A__ call_function getpathname strftime i2hex lldiv fwrite __window vfscanf rewind freopen njDecodeBlock pipe_read exit njUpsampleH pipe_r njGetImageSize __block_r atoi njGetImage __heap_r assert_fn gmtime strspn ctr0 drawstring_trans strlen __code toupper wcl njDone filename_cmp clock read_super_block abs strchr fputs acos strchrnul frexp vfprintf strpbrk read_sector free setpath njConvert  .symtab .strtab .shstrtab .text .data .got .got.plt .bss .eh_frame .comment                                                                                       �                                       !                �                                          '              @ �    @     `                              ,             `@ �   `@                                  5             �@ �   x@     �	                             :              P
 �    P      0                             D      0                �     *                                                   0�     @,      	   �                 	                      p�     u                                                   �     M                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      print("Hello, World!")
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         